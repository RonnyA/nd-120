/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : T_FLIPFLOP                                                   **
 **                                                                          **
 *****************************************************************************/

module T_FLIPFLOP( clock,
                   preset,
                   q,
                   qBar,
                   reset,
                   t,
                   tick );

   /*******************************************************************************
   ** Here all module parameters are defined with a dummy value                  **
   *******************************************************************************/
   parameter invertClockEnable = 1;

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input clock;
   input preset;
   input reset;
   input t;
   input tick;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output q;
   output qBar;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire s_clock;
   wire s_nextState;

   /*******************************************************************************
   ** The registers are defined here                                             **
   *******************************************************************************/
   reg s_currentState;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here the output signals are defined                                        **
   *******************************************************************************/
   assign q        = s_currentState;
   assign qBar     = ~(s_currentState);
   assign s_clock  = (invertClockEnable == 0) ? clock : ~clock;

   /*******************************************************************************
   ** Here the initial register value is defined; for simulation only            **
   *******************************************************************************/
   initial
   begin
      s_currentState = 0;
   end

   /*******************************************************************************
   ** Here the update logic is defined                                           **
   *******************************************************************************/
   assign s_nextState = s_currentState^t;

   /*******************************************************************************
   ** Here the actual state register is defined                                  **
   *******************************************************************************/
   //always @(posedge reset or posedge preset or posedge s_clock) //Vivado doesnt like ASYNC RESET )
   always @(posedge s_clock) //Vivado doesnt like ASYNC RESET )
   begin
      if (preset) s_currentState <= 1'b1;  // priority to pre-set
      else if (reset) s_currentState <= 1'b0;      
      else if (tick) s_currentState <= s_nextState;
   end

endmodule
