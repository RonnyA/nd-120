/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : F091                                                         **
 **                                                                          **
 *****************************************************************************/

module F091( N01,
             N02 );

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output N01;
   output N02;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire s_logisimNet0;
   wire s_logisimNet1;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign N01 = s_logisimNet0;
   assign N02 = s_logisimNet1;

   /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

   // Power
   assign  s_logisimNet0  =  1'b1;


   // Ground
   assign  s_logisimNet1  =  1'b0;


endmodule
