/**************************************************************************
** ND120 Shared                                                          **
**                                                                       **
** Component : MUX21L                                                    **
**                                                                       **
** Last reviewed: 11-NOV-2024                                            **
** Ronny Hansen                                                          **
***************************************************************************/

module MUX21L (
    input A,
    input B,
    input S,

    output ZN
);

  /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
  wire s_z;
  wire s_s;
  wire s_zn_out;
  wire s_a;
  wire s_b;

  /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

  /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
  assign s_s = S;
  assign s_a = A;
  assign s_b = B;

  /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
  assign ZN = s_zn_out;

  /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

  // NOT Gate
  assign s_zn_out = ~s_z;

  /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
  Multiplexer_2 PLEXERS_1 (
      .muxIn_0(s_a),
      .muxIn_1(s_b),
      .muxOut(s_z),
      .sel(s_s)
  );


endmodule
