/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : CPU_CS_PROM_19                                               **
 **                                                                          **
 *****************************************************************************/

module CPU_CS_PROM_19_ORG( input BLCS_n,         // Set to 0 to enable the output to IDB
                       input [1:0]  RF_1_0,  // Selects which of the 4 16 bit's of the microcoe to fetch
                       input [12:0] LUA_12_0, // Address of the microcode to fetch
                       
                       output [15:0] IDB_15_0 // The 16 bit microcode word
                       );


   wire [14:0] s_Address;
   wire [15:0] s_databus;

   assign s_Address[14:2] = LUA_12_0;
   assign s_Address[1:0]  = RF_1_0;


   // Controlled Buffer
   assign IDB_15_0 = (BLCS_n) ? 16'bZ : s_databus;


   // ROM: CHIP_23B_45132
   reg[7:0] s_CHIP_23B_45132_reg;
      always @(*)
      begin
         case (s_Address)
         {3'b000, 12'h000} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h001} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b000, 12'h002} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b000, 12'h004} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h006} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h008} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h00A} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h00C} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h00D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h00E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h00F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h010} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b000, 12'h011} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h012} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h013} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h014} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b000, 12'h015} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h016} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h017} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h018} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'h01A} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h01C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'h01E} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h020} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h022} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h024} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h026} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h028} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'h02A} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h02C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'h02E} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h030} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'h032} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h034} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h036} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h038} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b000, 12'h039} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h03A} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b000, 12'h03C} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b000, 12'h03D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b000, 12'h03E} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b000, 12'h03F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h040} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'h041} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'h042} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h043} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h046} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h047} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h049} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h04A} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h04E} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h051} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b000, 12'h052} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h053} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h055} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h056} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h058} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'h05A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h05B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h05C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h05D} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h05E} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h060} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b000, 12'h061} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b000, 12'h062} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b000, 12'h064} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h065} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h069} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h06B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h074} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h075} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h076} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h077} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h078} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b000, 12'h079} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h07A} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h07C} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b000, 12'h080} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'h081} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h084} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h085} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b000, 12'h086} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h087} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h088} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b000, 12'h089} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b000, 12'h08A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h08B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h08C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b000, 12'h08D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h090} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b000, 12'h094} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'h095} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h098} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'h099} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h09B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h09D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h09E} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h0A7} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h0A8} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b000, 12'h0AB} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h0AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h0AE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h0B7} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h0B8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h0BB} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h0BC} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b000, 12'h0BD} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h0BE} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h0BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0C2} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h0C5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h0C6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h0C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h0CA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h0CB} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b000, 12'h0CC} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b000, 12'h0CD} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h0CE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h0D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0D5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h0D6} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'h0D8} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b000, 12'h0D9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h0DA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h0DB} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'h0DC} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b000, 12'h0DD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h0DE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h0DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0E1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h0E2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0E4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b000, 12'h0E5} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h0E6} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h0E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0E9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h0EA} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h0EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0F2} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'h0F4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h0F5} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h0F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h0F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b000, 12'h0FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b000, 12'h100} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h104} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h106} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b000, 12'h108} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h10A} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h10C} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b000, 12'h10E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b000, 12'h110} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b000, 12'h112} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h114} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b000, 12'h115} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h116} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h118} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b000, 12'h119} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h11A} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h11C} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b000, 12'h11E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b000, 12'h120} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b000, 12'h122} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h124} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b000, 12'h125} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h126} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h128} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b000, 12'h129} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h12A} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h12C} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b000, 12'h12D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h12E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h130} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b000, 12'h131} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h132} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h134} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b000, 12'h135} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h136} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h138} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b000, 12'h139} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h13A} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h13C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b000, 12'h13D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h13E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h140} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b000, 12'h141} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h142} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h144} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b000, 12'h145} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h146} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h148} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b000, 12'h149} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h14A} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h14C} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b000, 12'h14D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h14E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h150} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b000, 12'h151} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h152} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h154} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h155} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h156} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h158} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h159} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h15A} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h15C} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'h15D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h15E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h160} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'h161} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h162} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h164} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b000, 12'h165} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h166} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h168} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b000, 12'h169} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h16A} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h16C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b000, 12'h16D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h16E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h170} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b000, 12'h171} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h172} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h174} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h175} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h176} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h178} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h179} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h17A} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h17C} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h17D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h17E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h180} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h181} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h182} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h184} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h185} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h186} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h188} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h189} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h18A} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h18D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h18E} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b000, 12'h191} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h192} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b000, 12'h195} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h196} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h198} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h19A} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h19C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h19E} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h1A0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h1A2} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h1A4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h1A6} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h1A8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h1AA} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h1AC} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b000, 12'h1AE} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h1B1} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h1B2} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b000, 12'h1B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h1B5} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b000, 12'h1B6} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h1B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h1B8} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b000, 12'h1B9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h1BA} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h1BC} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b000, 12'h1BE} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h1C0} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b000, 12'h1C2} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h1C4} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b000, 12'h1C5} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'h1C6} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b000, 12'h1C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h1C8} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b000, 12'h1C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h1CA} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h1CD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h1CE} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h1CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h1D1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h1D2} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h1D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h1D5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h1D6} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b000, 12'h1D9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h1DA} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b000, 12'h1DC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b000, 12'h1DD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h1DE} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h1E1} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h1E2} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h1E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h1E4} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b000, 12'h1E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h1E6} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h1E9} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'h1EA} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h1EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h1EC} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b000, 12'h1ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h1EE} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h1F1} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'h1F2} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h1F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h1F4} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b000, 12'h1F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h1F6} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h1F9} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h1FA} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h1FB} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h1FC} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b000, 12'h1FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h1FE} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h201} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h202} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h203} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h204} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h205} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h206} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h209} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h20A} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h20B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h20C} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'h20D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h20E} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h211} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h212} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h213} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h214} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b000, 12'h215} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h216} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h218} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b000, 12'h219} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h21A} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h21C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b000, 12'h21D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h21E} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b000, 12'h21F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h220} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h221} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b000, 12'h222} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b000, 12'h223} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h224} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h225} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b000, 12'h226} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b000, 12'h227} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h228} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h229} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h22A} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b000, 12'h22B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h22D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h22E} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b000, 12'h231} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h232} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h235} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h236} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b000, 12'h238} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h23A} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h23C} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h23E} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h244} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h248} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b000, 12'h24B} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b000, 12'h24C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h24D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h24E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b000, 12'h24F} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h250} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b000, 12'h253} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b000, 12'h254} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h255} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h256} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b000, 12'h257} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h258} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b000, 12'h259} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h25A} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b000, 12'h25C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h25D} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b000, 12'h25F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h260} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h265} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h268} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b000, 12'h269} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h26A} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b000, 12'h26C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h26D} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b000, 12'h26F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h270} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b000, 12'h271} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h272} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b000, 12'h274} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h275} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b000, 12'h277} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h278} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b000, 12'h279} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h27A} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b000, 12'h27D} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b000, 12'h27F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h280} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h281} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h284} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b000, 12'h285} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h287} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h288} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b000, 12'h289} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h28C} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b000, 12'h28D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h28E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h28F} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h290} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b000, 12'h293} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h294} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h296} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h29A} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h29B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h29C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h29F} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h2A0} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b000, 12'h2A1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h2A2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h2A3} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h2A4} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b000, 12'h2A7} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h2A8} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b000, 12'h2A9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h2AA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h2AB} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h2AC} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b000, 12'h2AF} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h2B0} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b000, 12'h2B1} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h2B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2B4} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b000, 12'h2B5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2BA} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h2BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2BC} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b000, 12'h2BF} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h2C0} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b000, 12'h2C1} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h2C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2C4} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b000, 12'h2C5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2CA} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h2CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2CF} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h2D0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h2D2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h2D3} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h2D4} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b000, 12'h2D5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2D9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h2DA} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h2DC} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b000, 12'h2DD} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h2DE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h2DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2E0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h2E1} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h2E3} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h2E5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h2E6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h2E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2EA} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h2EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2EC} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b000, 12'h2EF} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h2F0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h2F1} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h2F3} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h2F4} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b000, 12'h2F5} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h2F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2F8} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b000, 12'h2F9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h2FC} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b000, 12'h2FD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h2FE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h2FF} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h303} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h304} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b000, 12'h305} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h306} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h307} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h30B} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h30C} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b000, 12'h30D} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h30F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h310} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b000, 12'h311} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h315} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h316} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h318} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b000, 12'h319} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h31B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h31C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h31D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h320} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b000, 12'h321} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h322} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h323} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h324} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h327} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h328} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b000, 12'h329} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'h32A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h32B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h32C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h32F} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h330} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b000, 12'h331} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h333} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h334} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b000, 12'h335} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h339} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h33A} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h33C} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b000, 12'h33D} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h33F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h340} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h341} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h344} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b000, 12'h345} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h346} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h347} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h348} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h34B} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h34C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b000, 12'h34D} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'h34E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h34F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h350} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h353} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h354} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h355} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h357} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h358} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b000, 12'h35C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b000, 12'h35D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h362} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h363} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h368} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h36A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h36B} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h36C} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b000, 12'h36E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h370} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h371} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'h372} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h374} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h376} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h377} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h378} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b000, 12'h379} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h37A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h37B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h37C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h381} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h382} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h383} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'h389} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'h38A} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b000, 12'h38B} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h38D} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'h38E} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'h38F} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h391} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'h392} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'h393} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h395} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h396} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'h397} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h399} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b000, 12'h39A} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'h39B} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h39D} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b000, 12'h39E} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'h39F} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h3A2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h3A3} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3A6} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h3A8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h3A9} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b000, 12'h3AA} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'h3AB} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3AC} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h3B0} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h3B1} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'h3B2} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h3B5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h3B9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h3BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h3BE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'h3C0} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b000, 12'h3C1} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'h3C2} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b000, 12'h3C3} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3C4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b000, 12'h3C5} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'h3C6} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b000, 12'h3C7} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3C8} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b000, 12'h3C9} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'h3CA} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b000, 12'h3CB} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3CC} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b000, 12'h3CD} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h3CE} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b000, 12'h3CF} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3D0} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b000, 12'h3D1} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b000, 12'h3D2} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b000, 12'h3D3} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3D4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b000, 12'h3D5} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b000, 12'h3D6} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b000, 12'h3D7} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3D8} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b000, 12'h3D9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h3DA} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b000, 12'h3DB} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3DC} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b000, 12'h3DD} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b000, 12'h3DE} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b000, 12'h3DF} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3E0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h3E1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h3E4} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h3E9} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h3EA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h3EB} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'h3ED} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h3F0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h3F3} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h3F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h3F6} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b000, 12'h3F8} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h3FC} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h401} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h402} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h406} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h407} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h408} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b000, 12'h40A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h40B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h40C} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'h40D} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h40E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h40F} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'h410} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'h412} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h413} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h414} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h417} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h418} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'h41A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h41D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h41E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h41F} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h421} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h422} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h423} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b000, 12'h425} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h428} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h42C} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h431} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h432} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h435} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h438} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b000, 12'h43A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h43B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h43C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b000, 12'h43D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h440} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h443} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h445} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'h44B} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h450} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h451} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h452} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h453} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b000, 12'h454} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'h455} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h456} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h459} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h45A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h45B} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h45C} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b000, 12'h45F} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'h460} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b000, 12'h461} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h463} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b000, 12'h464} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'h465} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b000, 12'h468} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b000, 12'h469} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h46B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h46C} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b000, 12'h46D} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b000, 12'h46F} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b000, 12'h471} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h473} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h475} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h477} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h478} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b000, 12'h479} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h47B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h47C} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b000, 12'h47D} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b000, 12'h480} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h481} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b000, 12'h482} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b000, 12'h483} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h485} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h486} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h487} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h489} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h48A} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'h48B} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h48C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h48D} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h48E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'h48F} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h491} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b000, 12'h493} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h496} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h497} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h499} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h49C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h49D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h4A0} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h4A1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4A3} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h4A5} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h4A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4A8} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b000, 12'h4AC} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b000, 12'h4AD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4B0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b000, 12'h4B4} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h4B5} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b000, 12'h4B9} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h4BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4BC} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b000, 12'h4BD} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h4BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4C0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h4C1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4C5} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h4C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4C9} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h4CA} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h4CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h4CE} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h4CF} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h4D0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h4D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h4D3} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b000, 12'h4D4} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h4D6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4D8} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b000, 12'h4D9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4DA} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h4DB} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b000, 12'h4DD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h4DE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b000, 12'h4DF} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b000, 12'h4E1} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'h4E2} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b000, 12'h4E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4E4} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h4E5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h4E6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h4E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4E8} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b000, 12'h4E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h4EA} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h4ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h4EE} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h4F1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b000, 12'h4F2} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h4F4} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b000, 12'h4F9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h4FA} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h4FC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'h4FE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h4FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h501} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h504} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h505} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'h507} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h508} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h50A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h50C} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b000, 12'h50D} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b000, 12'h50F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h510} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h511} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h514} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b000, 12'h515} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h51E} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b000, 12'h521} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h522} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b000, 12'h523} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h524} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b000, 12'h525} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h526} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h527} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h528} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h529} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h52A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h52B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h52D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h52E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h531} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h532} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'h534} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b000, 12'h539} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h53E} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b000, 12'h53F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h540} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'h541} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h542} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h544} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h546} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h548} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b000, 12'h549} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b000, 12'h54A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h54E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h550} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h551} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b000, 12'h552} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h556} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h559} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b000, 12'h55B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h55D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h561} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h562} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h563} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h564} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h566} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h568} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b000, 12'h569} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h56A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h56C} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b000, 12'h56D} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b000, 12'h56E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h56F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h570} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b000, 12'h575} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h576} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h577} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h579} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h57B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h57C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h57E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h581} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'h582} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h583} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h585} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h587} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h588} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h58E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h590} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b000, 12'h591} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'h595} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h596} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h597} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h598} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'h599} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h59A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h59B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h59C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h5A1} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h5A2} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'h5A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5A4} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b000, 12'h5A5} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h5A6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5AA} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b000, 12'h5AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5AC} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b000, 12'h5AD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5B0} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b000, 12'h5B1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h5B2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5B4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h5B6} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b000, 12'h5B8} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b000, 12'h5B9} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b000, 12'h5BA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h5BC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b000, 12'h5BD} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h5BE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5C0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b000, 12'h5C4} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h5C5} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h5C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5C8} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b000, 12'h5C9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5CC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b000, 12'h5CD} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h5CE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5D0} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b000, 12'h5D2} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h5D5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h5D6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h5D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5D8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h5D9} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h5DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5DC} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b000, 12'h5DD} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'h5DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5E1} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h5E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5E4} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h5E5} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'h5E6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5E9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h5EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5EC} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b000, 12'h5EE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5F0} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b000, 12'h5F4} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h5F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h5F6} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h5F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5F8} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5F9} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b000, 12'h5FA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h5FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h5FD} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h5FE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h5FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h600} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h602} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h604} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b000, 12'h605} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'h606} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h607} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h608} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h609} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h60B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h60C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b000, 12'h60D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h60E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h610} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b000, 12'h611} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h615} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h616} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'h618} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b000, 12'h61A} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b000, 12'h61C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h61D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h61F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h620} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'h621} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'h622} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h623} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h625} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h628} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h629} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h62B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h62C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b000, 12'h62D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h630} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b000, 12'h631} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h634} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h638} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b000, 12'h63A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h63B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h63C} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b000, 12'h63D} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b000, 12'h640} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b000, 12'h641} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b000, 12'h644} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b000, 12'h645} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h648} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'h64C} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h650} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b000, 12'h652} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h653} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h654} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b000, 12'h655} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b000, 12'h658} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b000, 12'h659} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b000, 12'h65C} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b000, 12'h65D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h660} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'h664} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h665} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h669} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h676} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h677} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h678} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h67B} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h67C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b000, 12'h67D} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'h67E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h67F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h680} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b000, 12'h685} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h686} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h688} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b000, 12'h689} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b000, 12'h68A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h68B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h68C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b000, 12'h691} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h692} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h696} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h697} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h698} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h69B} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h69C} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b000, 12'h69D} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'h69E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h69F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h6A0} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h6A4} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b000, 12'h6A5} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b000, 12'h6A6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h6A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h6A8} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b000, 12'h6AD} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'h6AE} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b000, 12'h6B0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h6B4} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h6B8} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'h6BC} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h6C0} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h6C2} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h6C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h6C6} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h6C8} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b000, 12'h6C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h6CA} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h6CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h6CE} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h6D4} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b000, 12'h6D6} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h6D9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h6DA} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h6E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h6E2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'h6E5} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'h6E6} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h6E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h6EC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h6EE} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'h6F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h6F2} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h6F4} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h6F8} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b000, 12'h700} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h704} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b000, 12'h708} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h709} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h70A} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b000, 12'h70B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h70D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h70E} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h711} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h712} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b000, 12'h713} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h715} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h716} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h717} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h719} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h71A} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b000, 12'h71B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h71C} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b000, 12'h71D} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h71E} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'h722} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h723} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h725} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h726} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h729} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'h72A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h72B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h72C} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b000, 12'h72D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h72E} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h72F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h730} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b000, 12'h731} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'h732} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h733} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h736} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h738} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h739} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h73A} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h73C} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h73D} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b000, 12'h73E} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h73F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h741} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'h742} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h745} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h746} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h747} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h748} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h74A} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h74B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h74C} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b000, 12'h74D} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b000, 12'h74E} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h74F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h750} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b000, 12'h752} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h755} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b000, 12'h756} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b000, 12'h757} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h759} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h75A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h75B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h75C} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b000, 12'h75E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h762} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h764} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b000, 12'h766} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h767} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h768} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h769} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'h76A} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h76B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h76C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b000, 12'h76D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h76E} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h770} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b000, 12'h774} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b000, 12'h775} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h776} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h778} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b000, 12'h77C} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h77E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h782} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h788} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b000, 12'h789} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h78A} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h78B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h78C} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b000, 12'h78E} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h78F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h790} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b000, 12'h791} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'h792} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h793} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h795} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h79A} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b000, 12'h79D} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'h79E} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b000, 12'h79F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h7A0} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'h7A1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h7A2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h7AB} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h7AC} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b000, 12'h7AF} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h7B1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h7B6} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b000, 12'h7B8} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b000, 12'h7B9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h7BA} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h7BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h7BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h7BE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h7BF} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b000, 12'h7C1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h7C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h7C6} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h7C8} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b000, 12'h7C9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h7CA} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h7CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h7CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h7CE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h7CF} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'h7D0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h7D1} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h7D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h7D6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h7D8} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b000, 12'h7D9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h7DC} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b000, 12'h7DD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h7DE} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'h7E1} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'h7E2} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h7E4} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h7E5} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h7E9} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b000, 12'h7EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h7ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h7EE} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h7F5} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h7FA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h7FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h7FC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h7FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h7FE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h7FF} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'h801} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h805} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h806} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h808} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h80C} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h810} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'h814} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h815} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'h817} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h818} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b000, 12'h81A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h81D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h81E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h821} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h822} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b000, 12'h823} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h825} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b000, 12'h826} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h827} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h828} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h82A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h82C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h82D} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b000, 12'h82F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h830} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h831} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h832} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h833} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h835} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h837} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h839} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h83D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h83E} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h83F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h841} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h842} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h844} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b000, 12'h846} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h847} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h849} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h84C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h84D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h84E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h84F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h855} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h856} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h859} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h85C} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b000, 12'h85D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h85E} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h85F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h860} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b000, 12'h862} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h863} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h864} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h866} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h867} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h868} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b000, 12'h869} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h86C} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b000, 12'h86E} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h871} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h872} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h874} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h875} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h876} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h878} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'h879} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h87E} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b000, 12'h882} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b000, 12'h886} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b000, 12'h888} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b000, 12'h889} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h88A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h88B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h88C} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b000, 12'h88D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h88E} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b000, 12'h896} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'h89A} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'h89C} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'h89E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8A1} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'h8A2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h8A4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b000, 12'h8A5} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b000, 12'h8A6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h8A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8A8} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'h8AA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8AD} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b000, 12'h8AE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h8B0} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b000, 12'h8B1} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'h8B2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h8B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8B4} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b000, 12'h8B8} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b000, 12'h8B9} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b000, 12'h8BA} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'h8BC} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b000, 12'h8BD} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h8BE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h8BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8C4} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b000, 12'h8C5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h8C9} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h8CA} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'h8CC} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b000, 12'h8CD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h8D0} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'h8D2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8D4} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h8D5} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b000, 12'h8D6} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'h8D9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h8DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h8DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8DD} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h8DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'h8DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8E0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'h8E1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h8E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8E4} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b000, 12'h8E5} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b000, 12'h8E6} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b000, 12'h8E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8E8} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b000, 12'h8EC} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b000, 12'h8EE} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h8EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8F0} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'h8F1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8F2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h8F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h8F4} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b000, 12'h8F5} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h8F9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h8FA} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h8FD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b000, 12'h8FE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h901} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'h902} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h903} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h906} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h907} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h908} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h909} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'h90B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h90C} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b000, 12'h90D} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b000, 12'h90E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h910} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h911} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h913} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h914} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b000, 12'h915} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h916} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h918} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'h919} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'h91C} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b000, 12'h91D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h91E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h91F} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b000, 12'h922} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h923} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h926} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h92C} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b000, 12'h92D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'h92E} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h931} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'h932} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b000, 12'h933} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h934} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b000, 12'h935} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h936} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h937} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h938} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h939} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b000, 12'h93A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h93C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'h93D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h93E} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b000, 12'h93F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h941} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b000, 12'h943} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h944} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b000, 12'h947} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b000, 12'h94A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h94B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h94C} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b000, 12'h94E} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h950} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h951} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'h952} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'h953} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h956} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'h95C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b000, 12'h95E} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b000, 12'h961} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h962} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h964} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b000, 12'h965} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'h967} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h969} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h96A} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'h96C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h96D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h96E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'h970} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h971} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'h972} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h973} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h976} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h977} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b000, 12'h979} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'h97A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h97D} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'h97E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h97F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h982} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h983} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b000, 12'h984} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b000, 12'h986} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h987} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b000, 12'h989} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h98A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h98C} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b000, 12'h98E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h98F} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b000, 12'h990} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b000, 12'h991} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b000, 12'h992} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h993} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b000, 12'h995} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b000, 12'h996} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h997} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h999} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h99A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h99C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'h99D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h99E} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b000, 12'h9A0} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'h9A2} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'h9A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9A5} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h9A6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h9A7} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'h9AA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9AD} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b000, 12'h9AE} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'h9AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9B0} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'h9B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h9B2} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b000, 12'h9B5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b000, 12'h9B6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h9B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9B9} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h9BA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'h9BB} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'h9BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h9BE} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b000, 12'h9BF} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'h9C3} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h9C4} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b000, 12'h9C5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h9C6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9C9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h9CA} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h9CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9CC} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b000, 12'h9CE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9D0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'h9D2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h9D4} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'h9D5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9D6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h9D8} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b000, 12'h9DA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'h9DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9DD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9E0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b000, 12'h9E2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9E9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b000, 12'h9EA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'h9ED} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'h9EE} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'h9F1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'h9F4} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b000, 12'h9F5} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b000, 12'h9F6} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b000, 12'h9F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'h9F9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'h9FC} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b000, 12'h9FE} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'h9FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA01} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hA03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA04} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b000, 12'hA05} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b000, 12'hA06} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b000, 12'hA07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA08} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b000, 12'hA09} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'hA0A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hA0E} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'hA0F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA11} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hA13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA15} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hA16} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hA1A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hA1C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hA1E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hA20} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b000, 12'hA21} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'hA24} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b000, 12'hA25} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hA27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA28} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b000, 12'hA29} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hA2A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA2D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hA2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA31} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b000, 12'hA32} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hA34} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b000, 12'hA36} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hA37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA39} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hA3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA3C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b000, 12'hA3D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b000, 12'hA3E} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b000, 12'hA3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA40} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b000, 12'hA41} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'hA42} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hA43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA44} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b000, 12'hA45} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hA47} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA48} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b000, 12'hA49} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'hA4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA4C} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b000, 12'hA4D} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hA4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA55} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'hA56} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hA57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA59} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hA5A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hA5D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hA65} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hA66} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hA69} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hA6A} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b000, 12'hA6D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hA6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA71} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hA72} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hA73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA75} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hA79} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hA7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA7E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hA82} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hA83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA85} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hA87} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA89} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hA8A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hA8C} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b000, 12'hA8E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA8F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hA96} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hA9A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hA9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAA1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hAA2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hAA5} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hAA6} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hAA7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAAD} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hAAE} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hAAF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAB0} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b000, 12'hAB1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hAB2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAB3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAB5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hAB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAB9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hABA} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hABD} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hABE} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hABF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAC5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hAC6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hAC8} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b000, 12'hAC9} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hACA} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b000, 12'hACB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hACD} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b000, 12'hACE} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'hAD0} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hAD1} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hAD6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hAD7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAD9} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hADE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hADF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAE1} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hAE5} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hAE7} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hAE9} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'hAEB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAEC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hAED} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hAEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAF0} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b000, 12'hAF1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hAF6} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hAF8} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b000, 12'hAFA} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'hAFC} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b000, 12'hAFE} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hB00} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hB01} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hB03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB04} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b000, 12'hB05} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB09} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hB0A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hB0D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hB0E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hB0F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB10} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b000, 12'hB11} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hB12} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hB14} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'hB15} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hB17} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB18} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hB19} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB1E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hB20} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hB21} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB24} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hB25} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hB27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB28} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'hB29} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hB2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB2C} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'hB2D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB32} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hB34} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'hB35} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB38} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'hB39} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hB3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB3C} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'hB3D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hB3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB41} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hB43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB44} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hB45} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hB49} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hB4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB4D} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'hB4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB51} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hB53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB54} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'hB59} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hB5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB5C} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hB5D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hB61} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b000, 12'hB62} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hB63} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB65} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hB66} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hB67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB68} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b000, 12'hB69} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'hB6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB6D} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'hB6E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hB6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB70} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'hB72} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB74} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hB75} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'hB78} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b000, 12'hB79} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'hB7C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hB7D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hB7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB80} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b000, 12'hB81} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b000, 12'hB83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB85} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b000, 12'hB86} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b000, 12'hB88} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b000, 12'hB89} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hB8E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB8F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB91} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hB95} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b000, 12'hB96} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hB97} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hB98} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hB99} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hB9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB9C} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'hB9E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hB9F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBA1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'hBA3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBA4} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b000, 12'hBA5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hBA6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hBA8} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b000, 12'hBAC} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b000, 12'hBAD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hBB0} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hBB1} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b000, 12'hBB4} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b000, 12'hBB5} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'hBB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBB8} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hBB9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hBBB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBBC} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b000, 12'hBC1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hBC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBC5} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'hBC9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b000, 12'hBCA} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'hBCD} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hBCE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hBCF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBD1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hBD3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBD5} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hBD7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBD8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hBD9} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hBDB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBDC} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hBE1} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b000, 12'hBE2} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hBE3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBE6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hBE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBE8} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b000, 12'hBED} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hBEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBF0} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hBF4} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b000, 12'hBF5} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hBF7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBF8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hBF9} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hBFB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hBFD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hBFE} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hBFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC01} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hC02} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hC03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC04} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b000, 12'hC05} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hC07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC08} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hC0C} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b000, 12'hC0D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hC0F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC12} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hC13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC14} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'hC18} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b000, 12'hC19} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC1C} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b000, 12'hC24} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hC25} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hC26} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hC2A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC2D} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hC30} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'hC32} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC33} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC34} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hC35} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'hC39} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hC3A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hC3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC3D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hC3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC40} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b000, 12'hC41} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'hC45} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hC46} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hC47} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC49} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hC4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC4C} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hC4D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC50} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b000, 12'hC51} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hC53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC54} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b000, 12'hC55} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b000, 12'hC56} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hC59} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'hC5C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'hC5E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hC5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC60} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hC61} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b000, 12'hC63} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC65} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hC67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC69} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hC6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC6D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hC6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC71} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hC73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC76} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hC77} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC78} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hC79} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hC7A} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hC7C} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'hC7D} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b000, 12'hC7E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hC7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC81} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hC84} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b000, 12'hC85} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hC86} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hC87} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC88} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b000, 12'hC89} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hC8A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hC8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC8C} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hC8D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hC90} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hC91} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hC92} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hC93} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC94} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'hC95} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hC96} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hC97} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hC98} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hC9C} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hC9D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hCA0} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'hCA1} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hCA4} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hCA8} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b000, 12'hCAC} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b000, 12'hCAD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCB0} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b000, 12'hCB1} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b000, 12'hCB4} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b000, 12'hCB5} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'hCB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCB8} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b000, 12'hCB9} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b000, 12'hCBA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hCBB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCBC} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hCBD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hCBE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hCBF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCC1} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hCC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCC5} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'hCC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCC8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b000, 12'hCC9} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hCCB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCCC} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b000, 12'hCCD} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hCCF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCD0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b000, 12'hCD4} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b000, 12'hCD5} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hCD7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCD9} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b000, 12'hCDC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hCDD} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hCDF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCE1} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hCE3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCE4} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b000, 12'hCE5} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'hCE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCE8} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b000, 12'hCEC} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b000, 12'hCED} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hCEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCF0} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hCF1} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hCF5} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'hCF7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hCF8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hCF9} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hCFC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b000, 12'hCFD} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'hCFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD00} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b000, 12'hD01} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b000, 12'hD02} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hD03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD04} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b000, 12'hD08} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b000, 12'hD0C} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b000, 12'hD0D} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hD0F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD11} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b000, 12'hD14} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hD15} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hD17} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD19} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hD1B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD1C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b000, 12'hD1D} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'hD1F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD20} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b000, 12'hD21} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hD23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD24} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b000, 12'hD28} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b000, 12'hD2C} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b000, 12'hD30} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b000, 12'hD34} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hD35} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hD37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD38} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hD39} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b000, 12'hD3C} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b000, 12'hD3D} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'hD3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD40} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b000, 12'hD41} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b000, 12'hD42} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hD43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD44} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b000, 12'hD45} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hD47} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD48} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b000, 12'hD49} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hD4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD4C} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b000, 12'hD50} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b000, 12'hD51} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hD54} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hD55} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hD57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD58} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b000, 12'hD59} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD5C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hD5D} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hD5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD60} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b000, 12'hD61} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hD63} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD65} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b000, 12'hD68} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hD69} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hD6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD6D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hD6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD70} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b000, 12'hD71} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'hD73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD74} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b000, 12'hD78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b000, 12'hD79} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hD7D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b000, 12'hD80} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b000, 12'hD84} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b000, 12'hD85} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hD87} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD88} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b000, 12'hD89} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hD8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD8C} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b000, 12'hD90} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b000, 12'hD94} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b000, 12'hD95} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'hD97} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD98} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b000, 12'hD99} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b000, 12'hD9A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hD9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hD9C} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b000, 12'hDA0} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b000, 12'hDA4} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hDA5} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hDA7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDA8} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b000, 12'hDA9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDAC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hDAD} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hDAF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDB0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b000, 12'hDB1} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hDB3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDB5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDB8} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hDB9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hDBB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDBD} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hDBF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDC0} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b000, 12'hDC1} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'hDC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDC4} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b000, 12'hDC8} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b000, 12'hDCC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hDCD} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hDCF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDD0} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b000, 12'hDD2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hDD5} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hDD6} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'hDD7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDDA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hDDB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDDD} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b000, 12'hDDE} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b000, 12'hDE1} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b000, 12'hDE2} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hDE3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDE6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hDE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDEB} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hDEC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'hDED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hDEE} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'hDF1} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hDF2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hDF3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDF5} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hDF7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hDF8} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b000, 12'hDF9} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b000, 12'hDFA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hDFB} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hDFD} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b000, 12'hDFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE00} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b000, 12'hE01} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hE03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE04} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b000, 12'hE05} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hE07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE08} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hE09} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b000, 12'hE0A} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hE0B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE0C} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b000, 12'hE0D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE0E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hE10} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b000, 12'hE12} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hE13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE14} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b000, 12'hE15} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b000, 12'hE16} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hE17} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE19} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hE1A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hE1B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE1C} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b000, 12'hE20} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b000, 12'hE21} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE24} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b000, 12'hE25} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE29} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hE2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE2D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'hE31} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b000, 12'hE32} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hE34} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hE36} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hE37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE38} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b000, 12'hE39} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b000, 12'hE3C} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b000, 12'hE3D} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hE3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE41} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hE43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE45} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hE49} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hE4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE4C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hE4D} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b000, 12'hE4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE51} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hE52} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'hE54} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hE55} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hE56} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hE57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE58} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b000, 12'hE59} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hE5C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hE62} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hE64} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hE65} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE68} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'hE6A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE6D} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hE71} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hE73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE75} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hE77} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE78} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'hE79} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hE7A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE7C} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b000, 12'hE7D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hE7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE80} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'hE82} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE85} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hE8A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE8D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hE90} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b000, 12'hE91} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b000, 12'hE92} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b000, 12'hE95} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hE97} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hE99} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'hE9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE9C} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'hE9E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hE9F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEA1} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hEA5} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b000, 12'hEA6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hEA7} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hEA8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hEA9} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b000, 12'hEAB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEAC} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b000, 12'hEAD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEB1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hEB2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hEB5} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hEB6} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hEB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEB8} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b000, 12'hEB9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hEBA} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hEBC} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hEBD} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hEBF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEC0} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hEC1} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hEC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEC4} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b000, 12'hEC5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hEC8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hEC9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hECC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hED0} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'hED1} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'hED3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hED4} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hED5} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hED7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hED8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b000, 12'hED9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hEDB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEDC} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b000, 12'hEDD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hEE0} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hEE1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEE4} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hEE8} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'hEE9} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'hEEB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEEC} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hEED} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b000, 12'hEEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEF0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b000, 12'hEF1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hEF3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEF4} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hEF9} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hEFB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hEFE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hEFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF01} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hF03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF04} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b000, 12'hF05} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hF08} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hF09} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF0D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b000, 12'hF0E} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hF0F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF11} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b000, 12'hF12} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hF13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF14} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hF15} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hF18} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b000, 12'hF19} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b000, 12'hF1B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF1C} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b000, 12'hF1D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hF1F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF20} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b000, 12'hF21} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hF23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF24} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hF29} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hF2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF2E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hF2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF30} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b000, 12'hF31} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hF34} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b000, 12'hF35} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF39} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b000, 12'hF3A} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b000, 12'hF3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF3D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hF3E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b000, 12'hF3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF41} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hF43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF44} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b000, 12'hF45} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hF48} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b000, 12'hF49} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF4C} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b000, 12'hF4D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hF4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF50} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b000, 12'hF51} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hF53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF54} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'hF55} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'hF56} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'hF58} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hF5A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF5C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hF5D} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b000, 12'hF60} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'hF64} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b000, 12'hF65} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hF66} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b000, 12'hF67} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'hF68} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'hF6D} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hF6E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hF6F} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'hF70} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b000, 12'hF74} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b000, 12'hF75} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b000, 12'hF77} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF78} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hF79} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b000, 12'hF7A} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'hF7C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hF7D} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b000, 12'hF7E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hF7F} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hF81} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hF82} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b000, 12'hF83} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b000, 12'hF86} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hF87} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b000, 12'hF88} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hF89} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'hF8A} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'hF8C} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b000, 12'hF8D} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b000, 12'hF8E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b000, 12'hF8F} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b000, 12'hF91} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b000, 12'hF92} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b000, 12'hF93} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b000, 12'hF94} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b000, 12'hF95} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hF96} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b000, 12'hF97} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF98} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hF99} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b000, 12'hF9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hF9C} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b000, 12'hF9D} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b000, 12'hF9E} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b000, 12'hF9F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFA0} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b000, 12'hFA1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFA4} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'hFA5} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hFA6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hFA8} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'hFA9} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hFAA} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hFAC} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b000, 12'hFAD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFB0} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'hFB1} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b000, 12'hFB2} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hFB3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFB4} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b000, 12'hFB5} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b000, 12'hFB6} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hFB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFBC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b000, 12'hFBE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hFC1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFC5} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b000, 12'hFC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFC8} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b000, 12'hFCB} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b000, 12'hFCC} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b000, 12'hFCD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFD0} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFD5} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b000, 12'hFD6} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'hFD7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFD9} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b000, 12'hFDA} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'hFDB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFDD} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b000, 12'hFDE} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hFDF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFE5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b000, 12'hFE6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b000, 12'hFE9} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b000, 12'hFEA} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b000, 12'hFEB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFED} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b000, 12'hFEE} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b000, 12'hFEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFF1} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b000, 12'hFF2} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b000, 12'hFF3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b000, 12'hFF8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b000, 12'hFFA} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b000, 12'hFFC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b000, 12'hFFD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h000} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h001} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h003} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h004} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b001, 12'h005} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h006} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b001, 12'h007} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h008} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h009} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h00A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h00B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h00C} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b001, 12'h00D} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h00F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h012} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b001, 12'h013} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h016} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h01A} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h01D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h01E} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h020} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b001, 12'h022} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b001, 12'h026} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h027} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h029} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h02A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h02D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h02E} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b001, 12'h02F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h031} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h035} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h036} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h039} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h03A} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h03C} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b001, 12'h042} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b001, 12'h046} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'h048} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b001, 12'h04A} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b001, 12'h04E} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b001, 12'h052} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'h054} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'h056} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b001, 12'h058} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h060} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b001, 12'h061} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'h062} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h064} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b001, 12'h066} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h067} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h069} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h06A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h06D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h06E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h070} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b001, 12'h071} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h072} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'h07A} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h07D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h07E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h081} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h082} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h084} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b001, 12'h085} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h086} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h089} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h08A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h08D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h090} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b001, 12'h091} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h092} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b001, 12'h093} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h094} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b001, 12'h099} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b001, 12'h09A} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b001, 12'h09C} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b001, 12'h09D} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h09E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h0A0} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b001, 12'h0A1} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h0A2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h0A4} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b001, 12'h0A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h0A6} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b001, 12'h0A8} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h0AA} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h0AD} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h0AE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0B1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h0B5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h0B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0B8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h0B9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h0BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0BC} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h0BD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0C1} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h0C2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0C4} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h0C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h0C6} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'h0C8} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h0CD} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'h0D0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h0D1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h0D4} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h0D5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0D9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h0DA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0DC} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h0DD} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b001, 12'h0DE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h0E0} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b001, 12'h0E2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0E4} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b001, 12'h0E5} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'h0E6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0E9} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b001, 12'h0EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0EC} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b001, 12'h0EE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0F0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h0F4} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h0F5} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'h0F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0F8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h0FA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h0FC} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b001, 12'h0FD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h101} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h102} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h103} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h104} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b001, 12'h105} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h106} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h107} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h10B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h10C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h110} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h111} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b001, 12'h113} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h114} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b001, 12'h115} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h119} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h11A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h11B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h11E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h120} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h122} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h123} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h126} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h128} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h129} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h12D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h12E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h12F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h130} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h131} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h132} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'h135} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h136} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'h137} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h13C} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b001, 12'h13E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h13F} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'h140} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h141} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h142} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'h144} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b001, 12'h145} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'h147} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h148} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h14D} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'h14E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'h151} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h152} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'h153} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h155} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h156} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h157} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h158} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b001, 12'h159} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h15A} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'h15C} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b001, 12'h15D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h15E} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h15F} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'h160} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h162} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'h163} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h166} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h168} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h169} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b001, 12'h16A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h16B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h16C} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b001, 12'h16D} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b001, 12'h16E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h171} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h172} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h173} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h174} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b001, 12'h175} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h176} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h177} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h179} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h17A} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h17B} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'h17D} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h181} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h182} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h183} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h184} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b001, 12'h189} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h18A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h18C} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b001, 12'h190} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h192} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h194} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b001, 12'h19A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h19C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h1A0} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h1A1} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b001, 12'h1A2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h1A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1A4} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b001, 12'h1A5} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'h1A8} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'h1A9} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h1AC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b001, 12'h1AE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1B1} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h1B2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1B5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h1B6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1B8} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b001, 12'h1B9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h1BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h1BE} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h1C0} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'h1C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h1C2} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b001, 12'h1C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1C5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h1C6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1C9} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h1CA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1CC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b001, 12'h1CE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h1D1} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h1D2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1D5} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h1D6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1D9} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h1DA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1DC} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b001, 12'h1DD} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h1DE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h1E2} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h1E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h1E6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1E7} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'h1E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h1EA} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b001, 12'h1ED} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h1EE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1F1} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h1F2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1F5} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h1F6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1F9} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h1FA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h1FD} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h1FE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h201} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h202} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h205} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h206} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h208} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b001, 12'h209} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h20A} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'h20D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h20E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h210} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h211} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h212} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h213} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h214} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b001, 12'h215} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h216} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'h217} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h218} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h21A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h21C} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b001, 12'h21D} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b001, 12'h21E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h221} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h222} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b001, 12'h22B} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'h22C} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'h22F} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'h230} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h232} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h234} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h235} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h236} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h238} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b001, 12'h239} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h23A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h23B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h23D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h23E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h241} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h244} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h245} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h248} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h249} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h24C} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h24D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h250} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h251} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h252} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h253} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h254} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h255} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h256} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h257} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h259} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h25A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h25B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h25C} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h25D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h25E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h25F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h260} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h261} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h262} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h263} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h264} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h265} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h267} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h268} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b001, 12'h269} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'h26A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h26B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h26D} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h26F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h270} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b001, 12'h271} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h274} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h275} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h276} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'h278} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b001, 12'h279} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h27A} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b001, 12'h27B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h27C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h27D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h27E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h280} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b001, 12'h281} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b001, 12'h282} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h283} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h285} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h286} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b001, 12'h289} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h28A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h28F} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'h290} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'h293} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'h294} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b001, 12'h298} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b001, 12'h299} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h29C} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b001, 12'h29D} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h29E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h29F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2A0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h2A1} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b001, 12'h2A2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h2A4} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b001, 12'h2A8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h2A9} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h2AA} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b001, 12'h2AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2AC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h2AD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2B0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b001, 12'h2B4} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h2B5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2B8} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h2BA} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'h2BC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h2BD} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h2BE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h2BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2C0} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h2C1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2C4} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b001, 12'h2C8} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b001, 12'h2C9} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h2CD} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h2D0} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b001, 12'h2D1} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h2D2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h2D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2D4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h2D5} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h2D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2D8} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b001, 12'h2D9} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b001, 12'h2DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2DC} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b001, 12'h2DD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2E0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b001, 12'h2E5} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'h2E6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h2E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2E8} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b001, 12'h2E9} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h2EC} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b001, 12'h2ED} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b001, 12'h2F1} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h2F4} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b001, 12'h2F8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h2F9} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h2FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h2FC} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'h2FD} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b001, 12'h2FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h300} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b001, 12'h301} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b001, 12'h302} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'h303} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h304} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b001, 12'h308} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h309} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h30B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h30C} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h30D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h310} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b001, 12'h314} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h318} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h319} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h31C} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h31E} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'h320} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h321} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h322} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h323} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h324} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h325} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'h327} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h328} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b001, 12'h329} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h32C} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h32D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h330} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b001, 12'h331} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h332} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h333} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h334} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h335} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h336} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h337} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h338} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h339} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h33A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h33B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h33C} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b001, 12'h33D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h33E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h340} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b001, 12'h344} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b001, 12'h345} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h346} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h347} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h348} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b001, 12'h349} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h34A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'h34B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h34C} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b001, 12'h34E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h34F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h351} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'h354} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b001, 12'h355} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h357} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h358} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b001, 12'h359} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h35C} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b001, 12'h362} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'h364} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b001, 12'h366} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h367} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h36A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'h36B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h36D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'h36E} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h36F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h370} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b001, 12'h371} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h372} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h374} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b001, 12'h375} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h377} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h378} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b001, 12'h379} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h37D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h37E} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b001, 12'h381} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h384} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h385} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h386} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h387} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h388} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b001, 12'h389} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h38A} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'h38B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h38C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h38E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h390} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b001, 12'h391} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h392} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h394} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h396} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b001, 12'h398} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h399} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h39C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h39D} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h39E} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b001, 12'h39F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3A0} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b001, 12'h3A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h3A2} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'h3A4} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b001, 12'h3A5} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h3A8} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b001, 12'h3A9} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b001, 12'h3AA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h3AC} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b001, 12'h3AD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h3AE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h3AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3B0} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b001, 12'h3B1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3B4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h3B8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b001, 12'h3B9} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b001, 12'h3BA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h3BD} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h3BE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h3BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3C1} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h3C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3C5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h3C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3C9} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h3CA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h3CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3CC} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b001, 12'h3CE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3D0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b001, 12'h3D2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3D4} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b001, 12'h3D5} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h3D6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h3D8} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b001, 12'h3DA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h3DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3DC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h3DD} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h3DE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h3DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3E0} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b001, 12'h3E1} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b001, 12'h3E2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h3E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3E4} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b001, 12'h3E5} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h3E8} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b001, 12'h3E9} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h3ED} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b001, 12'h3EE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h3EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3F0} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b001, 12'h3F1} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h3F2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h3F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3F4} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'h3F8} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b001, 12'h3F9} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h3FA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h3FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h3FC} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b001, 12'h3FD} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h3FE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h3FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h400} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h401} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h402} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h404} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'h405} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'h409} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h40A} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b001, 12'h40C} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b001, 12'h411} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h412} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h413} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h414} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b001, 12'h415} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h416} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h417} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h419} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h41A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h41B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h41C} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b001, 12'h41D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h41E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h420} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'h421} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h424} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h426} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h427} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h429} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h42A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h42C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b001, 12'h42D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h42E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h42F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h430} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'h431} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h434} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h435} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h437} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h438} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h439} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h43C} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h43E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h43F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h441} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h442} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h444} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b001, 12'h445} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h446} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h448} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b001, 12'h44A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h44D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h44E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h44F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h450} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b001, 12'h452} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h455} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h456} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'h457} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h458} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h45A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h45C} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h45D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h460} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h461} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h465} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h466} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h468} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'h469} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h46C} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b001, 12'h46E} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b001, 12'h472} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b001, 12'h473} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h474} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b001, 12'h476} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h47A} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b001, 12'h47C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h47D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h47E} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h480} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b001, 12'h481} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h485} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h487} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h488} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h489} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h48A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h48C} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b001, 12'h48D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h490} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b001, 12'h491} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h492} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h494} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b001, 12'h495} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h497} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h498} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b001, 12'h499} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h49C} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b001, 12'h49E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4A0} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h4A1} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b001, 12'h4A4} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b001, 12'h4A6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4A8} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b001, 12'h4A9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4AC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h4AE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h4B0} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'h4B1} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b001, 12'h4B4} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b001, 12'h4B5} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b001, 12'h4B8} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'h4B9} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b001, 12'h4BC} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b001, 12'h4BD} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'h4C0} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h4C1} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b001, 12'h4C4} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'h4C5} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'h4C6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4C8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h4C9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h4CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4CC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h4CD} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h4D0} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b001, 12'h4D1} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'h4D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4D4} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'h4D5} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h4D8} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b001, 12'h4D9} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h4DC} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b001, 12'h4DD} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h4E0} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b001, 12'h4E1} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'h4E4} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b001, 12'h4E5} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h4E8} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b001, 12'h4E9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4EC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h4EE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4F0} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h4F1} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h4F2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h4F4} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b001, 12'h4F5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4F8} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b001, 12'h4F9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h4FD} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h4FE} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b001, 12'h500} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b001, 12'h501} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h502} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h503} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h504} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h508} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h509} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'h50A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h50B} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b001, 12'h50C} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b001, 12'h50D} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b001, 12'h50E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h511} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h512} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b001, 12'h513} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h515} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'h516} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h518} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b001, 12'h519} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h51A} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h51B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h51C} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b001, 12'h51D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'h51E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h51F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h525} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h526} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'h528} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b001, 12'h52A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'h52B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h52D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h52E} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b001, 12'h530} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h531} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h532} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h533} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b001, 12'h535} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h537} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h539} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b001, 12'h53A} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b001, 12'h53B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h53C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h53D} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h53F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h540} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'h541} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'h542} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h543} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h545} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h546} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h549} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h54A} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h54D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h54E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h550} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h558} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b001, 12'h559} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h55D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h55E} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h561} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h562} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h568} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b001, 12'h569} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h56A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h56B} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b001, 12'h56D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h56E} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h571} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h572} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h574} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b001, 12'h578} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b001, 12'h57C} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b001, 12'h581} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h582} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h583} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h584} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b001, 12'h585} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h586} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h587} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h588} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b001, 12'h589} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h58A} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h58C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h58E} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h592} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h596} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b001, 12'h598} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b001, 12'h599} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h59A} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h59D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h5A1} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h5A2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h5A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5A4} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h5A6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5A8} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b001, 12'h5AA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5AD} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h5AE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h5B0} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h5B2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5B5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h5B6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h5B8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h5B9} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h5BA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h5BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5BC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h5BD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5C0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b001, 12'h5C4} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h5C5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5C9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'h5CA} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h5CC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h5CD} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h5CE} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b001, 12'h5D0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h5D1} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h5D2} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b001, 12'h5D4} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h5D5} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h5D6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h5D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5D9} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b001, 12'h5DA} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h5DD} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h5DE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h5DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5E1} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b001, 12'h5E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5E9} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h5EA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h5EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5ED} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h5EE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h5F0} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b001, 12'h5F1} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h5F2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h5F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5F5} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h5F6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h5F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5F9} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h5FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h5FD} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h5FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h601} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h603} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h604} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b001, 12'h605} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h606} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h607} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h60D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h60E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h611} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h612} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h613} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h615} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h616} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'h618} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b001, 12'h61C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h621} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h622} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h623} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h624} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b001, 12'h626} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h628} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'h629} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h62A} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'h62D} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h62E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h631} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h632} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h635} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h636} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h638} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b001, 12'h639} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h63A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h63C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h63D} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h63E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h640} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h641} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h642} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b001, 12'h644} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b001, 12'h645} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h646} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h647} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h648} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b001, 12'h64A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h64B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h64D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h651} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h653} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h654} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h655} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h656} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h657} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h658} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h659} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h65A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h65B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h65C} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h65D} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b001, 12'h65E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h65F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h660} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h661} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h662} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h663} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h664} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h665} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h666} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'h668} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'h669} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h66C} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b001, 12'h66D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h671} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h672} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b001, 12'h675} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h679} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h67A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h67B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h67D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h681} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h685} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h688} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h68C} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b001, 12'h68D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h690} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'h691} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h694} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b001, 12'h695} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b001, 12'h697} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h699} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h69B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h69C} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b001, 12'h69E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'h6A1} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h6A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h6A6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'h6A8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h6A9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h6AA} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b001, 12'h6AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6AC} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b001, 12'h6AD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6B0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h6B1} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b001, 12'h6B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6B4} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b001, 12'h6B5} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h6B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6B8} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h6B9} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h6BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6BD} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h6BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6C0} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b001, 12'h6C1} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h6C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6C4} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b001, 12'h6C5} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h6C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6C8} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b001, 12'h6C9} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'h6CA} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'h6CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6CC} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b001, 12'h6CD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6D0} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h6D1} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h6D2} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b001, 12'h6D5} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h6D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'h6D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6D9} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h6DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6DD} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h6DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6E0} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h6E1} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h6E5} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h6E6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h6E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6E9} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h6EA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h6EC} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'h6ED} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h6EE} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'h6F0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h6F1} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h6F2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h6F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h6F4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h6F5} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b001, 12'h6F6} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b001, 12'h6FA} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h6FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h6FE} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b001, 12'h700} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h701} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h702} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h703} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h704} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h705} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b001, 12'h706} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h707} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h708} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b001, 12'h709} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h70E} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'h712} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'h715} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h716} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b001, 12'h718} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'h719} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h71A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h71C} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b001, 12'h720} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b001, 12'h721} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h724} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h728} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h729} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h72A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h72B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h72C} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h72D} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b001, 12'h72E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h72F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h731} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h732} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h735} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h736} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h738} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h739} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h73A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h73C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b001, 12'h73D} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h73E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h73F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h740} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'h745} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h746} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h748} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b001, 12'h749} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h74A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h74B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h74C} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'h74D} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b001, 12'h74E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h74F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h750} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b001, 12'h752} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h754} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b001, 12'h755} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h756} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h758} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'h759} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h75B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h75D} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h75E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h761} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h762} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h764} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h766} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h767} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h769} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h76A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h76C} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b001, 12'h76D} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h76E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h771} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h774} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b001, 12'h775} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b001, 12'h778} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h779} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h77A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h77B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h77C} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b001, 12'h77D} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b001, 12'h77E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h77F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h781} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h784} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h785} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h786} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h788} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'h789} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h78A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h78B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h78D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h78F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h792} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h794} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b001, 12'h798} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h79A} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h79C} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b001, 12'h79D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7A1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h7A2} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h7A4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h7A5} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h7A6} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b001, 12'h7A8} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h7AC} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b001, 12'h7AE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7B0} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b001, 12'h7B1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7B4} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h7B8} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b001, 12'h7BA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7BC} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b001, 12'h7BD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7C0} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h7C2} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b001, 12'h7C4} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b001, 12'h7C6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7C8} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b001, 12'h7C9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7CC} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h7CE} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'h7D1} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h7D2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h7D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7D4} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b001, 12'h7D5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7D9} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h7DA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h7DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7DC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h7DD} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b001, 12'h7DE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h7DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7E0} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h7E1} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b001, 12'h7E2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h7E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7E4} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b001, 12'h7E5} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h7E6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h7E8} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b001, 12'h7EC} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'h7F0} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h7F2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7F4} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'h7F5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7F8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h7F9} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h7FA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h7FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h7FC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h7FD} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b001, 12'h7FE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h7FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h800} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h801} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h804} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b001, 12'h805} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h806} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b001, 12'h809} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h80A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h80B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h80C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b001, 12'h80D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h80E} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b001, 12'h810} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b001, 12'h814} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h815} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'h818} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b001, 12'h819} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h81A} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b001, 12'h81B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h81C} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h81D} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b001, 12'h81E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h81F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h820} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'h823} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h824} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h827} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'h828} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'h829} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h82A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h82B} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b001, 12'h82C} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h82D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h82E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h82F} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h830} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b001, 12'h832} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h834} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h837} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h838} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h839} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h83C} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b001, 12'h83D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h841} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h842} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h843} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h845} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'h846} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h849} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h84A} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h84D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h84E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h851} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h852} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h853} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h854} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h855} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h856} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h857} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b001, 12'h858} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'h859} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h85C} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h85D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h861} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h862} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b001, 12'h863} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h865} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h866} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h869} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h86A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h86B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h86C} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h86D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h870} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b001, 12'h871} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h872} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h875} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h876} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h877} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h878} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b001, 12'h879} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h87A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h87C} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'h87D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h880} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h881} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h882} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h883} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h884} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b001, 12'h885} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h886} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h888} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b001, 12'h88A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h88C} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h88D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h890} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h891} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h892} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h893} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h895} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h896} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h898} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h89A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h89B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h89D} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'h89E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h8A0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h8A1} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'h8A2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h8A5} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h8A6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h8A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h8A9} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h8AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h8AD} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h8AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h8B1} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h8B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h8B5} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h8B6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h8B9} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'h8BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h8BD} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h8BE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h8C1} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h8C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h8C4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h8C5} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h8C6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h8C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h8C8} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b001, 12'h8C9} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'h8CC} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b001, 12'h8CD} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'h8D0} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b001, 12'h8D1} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b001, 12'h8D4} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b001, 12'h8D5} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h8D8} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b001, 12'h8D9} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'h8DC} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b001, 12'h8DD} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b001, 12'h8E0} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b001, 12'h8E1} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'h8E4} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b001, 12'h8E5} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'h8E8} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b001, 12'h8E9} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'h8EC} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b001, 12'h8ED} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'h8F0} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b001, 12'h8F1} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'h8F4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'h8F5} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b001, 12'h8F8} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b001, 12'h8F9} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'h8FC} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b001, 12'h8FD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h8FE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h900} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b001, 12'h901} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h902} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h904} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b001, 12'h908} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b001, 12'h90B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h90C} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b001, 12'h90D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'h90F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h910} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b001, 12'h911} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'h913} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h914} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b001, 12'h915} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h917} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h918} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b001, 12'h919} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'h91B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h91C} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b001, 12'h91D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h91F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h920} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b001, 12'h921} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h923} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h924} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b001, 12'h925} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b001, 12'h927} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h928} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b001, 12'h929} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h92C} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b001, 12'h92D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h92E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h92F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h930} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b001, 12'h931} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h932} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h933} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h935} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h936} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h937} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h938} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b001, 12'h939} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h93A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h93B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h93D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h941} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h942} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h943} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h945} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h946} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h949} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h94A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h94D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h94E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h94F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h951} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h952} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h955} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h956} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h959} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h95A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h95C} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b001, 12'h95D} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'h95E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h960} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b001, 12'h961} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'h962} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h963} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h964} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b001, 12'h965} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'h966} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h968} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b001, 12'h969} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h96A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h96B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h96C} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b001, 12'h96D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h970} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'h975} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'h979} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h97A} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b001, 12'h97B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h97D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h981} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'h982} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h983} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h984} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b001, 12'h985} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h988} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b001, 12'h98C} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h98D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'h990} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b001, 12'h992} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h993} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h994} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b001, 12'h996} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h997} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h998} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b001, 12'h999} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'h99A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h99B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h99D} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h99F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9A0} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'h9A1} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'h9A2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'h9A4} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b001, 12'h9A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h9A6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h9A7} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b001, 12'h9AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h9AE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'h9B0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'h9B2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h9B4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b001, 12'h9B5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9B6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h9B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9B8} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'h9B9} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h9BA} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h9BD} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h9BE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9C1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h9C2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9C4} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b001, 12'h9C5} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'h9C6} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'h9C9} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h9CA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9CE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9D1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h9D2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9D4} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b001, 12'h9D5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9D9} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'h9DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b001, 12'h9E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b001, 12'h9E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b001, 12'h9E9} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b001, 12'h9EA} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'h9ED} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'h9EE} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'h9F1} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b001, 12'h9F2} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b001, 12'h9F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9F4} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'h9F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'h9F6} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'h9F8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'h9FA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'h9FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'h9FC} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b001, 12'h9FD} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b001, 12'h9FE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'h9FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA00} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b001, 12'hA01} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'hA02} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hA03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA04} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hA05} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hA08} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'hA09} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b001, 12'hA0A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hA0B} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hA0C} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b001, 12'hA0E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA0F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA10} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hA11} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA12} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA14} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b001, 12'hA15} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b001, 12'hA17} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA18} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'hA19} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hA1A} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hA1C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hA20} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b001, 12'hA21} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hA22} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hA24} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'hA25} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'hA26} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hA27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA29} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hA2A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA2D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hA2E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA30} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b001, 12'hA31} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hA32} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA33} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA34} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hA36} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hA38} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'hA39} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b001, 12'hA3A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hA3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA3D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hA3E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA41} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hA42} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA45} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hA48} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b001, 12'hA49} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hA4A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA4C} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'hA4D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'hA4E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hA4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA51} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hA52} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA55} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hA56} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA59} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hA5A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA5C} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA5D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hA5E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hA61} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hA62} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA63} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA64} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b001, 12'hA65} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hA66} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA68} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA69} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hA6A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hA6D} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hA6E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA70} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hA71} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hA72} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b001, 12'hA73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA75} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b001, 12'hA77} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hA79} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hA7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA7C} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b001, 12'hA7D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hA7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA80} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b001, 12'hA81} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'hA82} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hA83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA85} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hA87} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hA88} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hA89} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hA8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA8D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hA8F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA90} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b001, 12'hA91} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b001, 12'hA92} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hA95} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hA96} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA97} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA99} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hA9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hA9C} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hA9D} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b001, 12'hA9E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hAA5} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hAA6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hAA7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hAA8} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b001, 12'hAA9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hAAA} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hAAC} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hAB1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hAB2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hAB3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hAB4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hAB5} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hAB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hAB9} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hABC} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hABD} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hAC1} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hAC3} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hAC4} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b001, 12'hAC5} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hAC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hAC8} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b001, 12'hAC9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hACD} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hACF} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hAD0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b001, 12'hAD1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hAD5} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hAD6} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hAD9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hADA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hADB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hADD} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hADF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hAE0} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b001, 12'hAE1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'hAE2} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hAE3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hAE4} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hAE5} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hAE6} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hAE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hAE8} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b001, 12'hAE9} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'hAEB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hAEC} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b001, 12'hAED} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b001, 12'hAF1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hAF4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hAF5} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hAF8} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b001, 12'hAF9} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hAFA} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'hAFB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hAFD} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b001, 12'hAFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB01} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hB03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB05} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hB07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB08} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hB0B} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'hB0C} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hB0D} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'hB0E} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hB11} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hB13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB15} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b001, 12'hB17} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB18} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'hB19} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hB1A} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hB1D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hB21} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b001, 12'hB22} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hB23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB25} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hB26} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hB27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB28} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b001, 12'hB29} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hB2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB2C} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hB32} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hB33} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB34} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b001, 12'hB35} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'hB37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB38} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hB39} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hB3A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hB3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB3D} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b001, 12'hB3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB41} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hB44} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hB47} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'hB48} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hB49} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'hB4A} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hB4D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hB4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB51} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b001, 12'hB53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB54} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b001, 12'hB55} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b001, 12'hB56} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hB59} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hB5A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hB5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB5C} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hB5D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hB5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB61} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'hB62} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b001, 12'hB63} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB65} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'hB66} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hB67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB68} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'hB69} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'hB6A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hB6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB6C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hB6E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hB6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB70} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b001, 12'hB71} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'hB72} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hB73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB75} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hB76} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hB77} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB78} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b001, 12'hB79} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB7D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hB7E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB80} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b001, 12'hB81} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hB83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB84} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b001, 12'hB85} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b001, 12'hB86} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hB87} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB89} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hB8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB8D} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hB8E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hB8F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB90} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hB94} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b001, 12'hB95} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b001, 12'hB96} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hB97} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hB99} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hB9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBA0} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b001, 12'hBA1} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'hBA2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hBA3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBA5} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hBA7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBA9} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hBAB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBAD} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'hBAF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBB1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hBB2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hBB3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBB5} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'hBB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBB9} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hBBB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBBC} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hBC0} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hBC1} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'hBC2} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hBC7} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hBC9} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b001, 12'hBCB} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hBCD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hBCE} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hBD1} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hBD2} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hBD7} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hBD9} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b001, 12'hBDB} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hBDF} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hBE0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hBE1} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hBE3} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hBE5} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'hBE6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hBE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBE9} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'hBEB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBEC} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hBED} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b001, 12'hBF0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hBF4} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b001, 12'hBF5} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'hBF9} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hBFB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hBFC} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b001, 12'hBFD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hBFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC00} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hC05} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hC07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC09} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hC0B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC0D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hC10} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hC11} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hC13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC15} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'hC16} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b001, 12'hC17} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC19} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'hC1A} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hC1B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC1D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'hC20} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b001, 12'hC21} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hC22} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hC24} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hC26} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hC27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC28} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b001, 12'hC29} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b001, 12'hC2A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hC2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC2D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hC2E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hC2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC30} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b001, 12'hC35} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hC37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC38} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hC39} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC3A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hC3E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hC41} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hC42} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC44} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hC48} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b001, 12'hC49} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'hC4A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hC4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC4C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hC4D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hC4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC50} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b001, 12'hC51} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'hC53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC54} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hC58} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b001, 12'hC59} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b001, 12'hC5A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hC5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC5C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hC5D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hC5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC60} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b001, 12'hC61} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC64} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b001, 12'hC68} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hC69} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hC6A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC6D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'hC6E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hC6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC71} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hC72} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hC73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC74} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'hC75} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'hC76} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hC77} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC79} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hC7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC7D} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b001, 12'hC7E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hC7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC80} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hC81} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hC82} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hC83} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hC87} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hC89} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hC8B} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hC8F} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hC91} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b001, 12'hC93} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hC95} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hC96} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hC97} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hC98} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hC99} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hC9A} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hC9F} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hCA1} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b001, 12'hCA3} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hCA4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hCA5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hCA7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCA8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b001, 12'hCA9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCAA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hCAB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCAD} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hCAF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCB1} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b001, 12'hCB2} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hCB6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hCB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCB9} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hCBA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hCBB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCBC} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b001, 12'hCBD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hCBE} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hCC1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hCC2} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hCC4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hCC7} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hCC9} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b001, 12'hCCA} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hCCD} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hCCE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hCCF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCD0} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hCD1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hCD3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCD5} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hCD8} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b001, 12'hCD9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hCDA} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hCDD} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hCDE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hCDF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCE0} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'hCE2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCE3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCE4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hCE5} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b001, 12'hCE8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hCE9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hCED} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hCEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCF0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b001, 12'hCF1} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b001, 12'hCF5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hCF8} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b001, 12'hCF9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hCFB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hCFD} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hCFE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hCFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD00} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b001, 12'hD01} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b001, 12'hD06} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hD07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD08} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hD0C} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b001, 12'hD0D} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'hD11} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hD12} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b001, 12'hD15} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hD16} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hD18} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b001, 12'hD1C} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b001, 12'hD1D} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hD1E} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hD21} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hD22} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hD23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD25} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hD27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD28} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b001, 12'hD29} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'hD2A} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hD2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD2D} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b001, 12'hD2F} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hD31} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hD33} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD37} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'hD38} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'hD39} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'hD3A} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hD3C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hD3D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hD3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD41} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b001, 12'hD43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD45} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hD49} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hD4A} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b001, 12'hD4C} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'hD4D} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b001, 12'hD4E} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b001, 12'hD4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD50} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hD51} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hD52} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hD53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD55} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b001, 12'hD57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD59} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b001, 12'hD5A} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hD5D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hD5E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hD5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD61} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hD63} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD64} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hD65} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hD66} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD69} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hD6A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD6C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hD6D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hD6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD70} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b001, 12'hD71} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hD72} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hD74} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hD76} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hD78} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b001, 12'hD79} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD7C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hD7D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hD7E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hD7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD81} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b001, 12'hD83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD85} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hD87} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD88} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hD89} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hD8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD8C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hD8D} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b001, 12'hD8F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD91} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hD93} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hD95} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hD99} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b001, 12'hD9A} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b001, 12'hD9C} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b001, 12'hD9D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hDA0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b001, 12'hDA4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b001, 12'hDA8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b001, 12'hDAC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b001, 12'hDB0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b001, 12'hDB4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b001, 12'hDB8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b001, 12'hDBC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b001, 12'hDC2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDC4} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'hDC6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDC8} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hDCA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDCB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDCC} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hDCE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDCF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDD2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDD3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDD4} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDD6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDD7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDD8} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'hDDA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDDB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDDE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDDF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDE2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDE3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDE4} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'hDE6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDE8} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hDEA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDEB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDEC} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hDEE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDF2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDF3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDF4} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDF6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDF7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDF8} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b001, 12'hDFA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDFB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDFE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hDFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hE00} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b001, 12'hE01} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE02} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'hE04} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b001, 12'hE05} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE06} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'hE08} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b001, 12'hE09} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE0A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'hE0C} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b001, 12'hE0D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE0E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'hE10} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hE12} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'hE14} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hE16} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'hE18} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b001, 12'hE1A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'hE1C} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b001, 12'hE1E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'hE20} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b001, 12'hE21} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE22} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'hE24} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b001, 12'hE25} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE26} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'hE28} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b001, 12'hE29} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE2A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'hE2C} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b001, 12'hE2D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE2E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'hE30} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hE32} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'hE34} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hE36} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'hE38} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b001, 12'hE3A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'hE3C} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b001, 12'hE3E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'hE40} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b001, 12'hE44} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b001, 12'hE45} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hE46} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b001, 12'hE48} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b001, 12'hE49} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hE4A} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b001, 12'hE4C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b001, 12'hE4D} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hE50} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hE51} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'hE52} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b001, 12'hE53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hE54} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b001, 12'hE55} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b001, 12'hE56} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hE57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hE58} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b001, 12'hE59} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'hE5A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'hE5C} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b001, 12'hE5D} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b001, 12'hE5E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hE5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hE60} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hE64} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b001, 12'hE65} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hE66} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hE67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hE68} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b001, 12'hE69} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'hE6A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'hE6D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'hE6E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hE6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hE71} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b001, 12'hE72} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'hE74} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'hE75} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'hE76} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'hE78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b001, 12'hE7C} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hE7D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'hE7E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hE7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hE80} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b001, 12'hE84} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b001, 12'hE86} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE88} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b001, 12'hE8A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE8C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hE8E} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'hE90} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b001, 12'hE92} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE94} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b001, 12'hE96} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE98} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b001, 12'hE9A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hE9C} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b001, 12'hE9E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hEA0} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b001, 12'hEA2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hEA4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hEA6} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'hEA8} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b001, 12'hEAA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hEAC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hEAE} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'hEB0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hEB2} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'hEB4} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b001, 12'hEB8} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b001, 12'hEB9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hEBA} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hEBC} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b001, 12'hEBD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hEBE} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b001, 12'hEC1} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hEC2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hEC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hEC5} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hEC6} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b001, 12'hEC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hEC8} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b001, 12'hEC9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'hECA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hECB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hECC} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b001, 12'hECD} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'hECE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hECF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hED0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b001, 12'hED1} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'hED2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hED3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hED4} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b001, 12'hED5} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hED6} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b001, 12'hED7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hED8} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b001, 12'hED9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'hEDA} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b001, 12'hEDB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hEDC} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b001, 12'hEDD} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'hEDE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hEDF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hEE1} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hEE2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hEE3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hEE5} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hEE6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hEE7} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b001, 12'hEE8} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b001, 12'hEE9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hEEA} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b001, 12'hEEC} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b001, 12'hEED} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hEEE} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hEEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hEF0} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b001, 12'hEF4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b001, 12'hEF5} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hEF6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b001, 12'hEF7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hEF9} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hEFC} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b001, 12'hEFE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hEFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF00} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hF07} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b001, 12'hF08} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b001, 12'hF0C} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b001, 12'hF0E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hF10} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'hF14} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b001, 12'hF18} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b001, 12'hF19} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b001, 12'hF1A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'hF1C} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b001, 12'hF1D} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b001, 12'hF1E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b001, 12'hF20} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b001, 12'hF22} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hF23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF24} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b001, 12'hF28} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b001, 12'hF2D} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b001, 12'hF2E} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b001, 12'hF2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF30} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'hF34} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b001, 12'hF38} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b001, 12'hF3C} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hF3E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hF3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF40} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b001, 12'hF41} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hF42} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b001, 12'hF43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF48} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b001, 12'hF4A} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b001, 12'hF4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF4C} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b001, 12'hF4D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b001, 12'hF4E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hF4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF51} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hF56} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hF58} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b001, 12'hF59} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hF5C} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b001, 12'hF5D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b001, 12'hF5E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b001, 12'hF5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF64} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b001, 12'hF66} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hF68} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b001, 12'hF69} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b001, 12'hF6A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF6C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b001, 12'hF6E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b001, 12'hF70} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b001, 12'hF74} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b001, 12'hF78} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b001, 12'hF7C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b001, 12'hF80} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b001, 12'hF81} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b001, 12'hF83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF84} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b001, 12'hF85} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b001, 12'hF87} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF88} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b001, 12'hF89} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b001, 12'hF8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF8C} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b001, 12'hF8D} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hF8F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF90} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hF91} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hF93} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF94} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hF95} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hF97} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF98} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hF99} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hF9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hF9C} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hF9D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hF9F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFA0} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hFA1} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hFA3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFA4} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hFA5} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hFA7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFA8} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hFA9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hFAB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFAC} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hFAD} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hFAF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFB0} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hFB1} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hFB3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFB4} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hFB5} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hFB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFB8} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b001, 12'hFB9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b001, 12'hFBB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFBC} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b001, 12'hFBD} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b001, 12'hFBF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFC0} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'hFC1} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hFC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFC4} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b001, 12'hFC5} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hFC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFC8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b001, 12'hFC9} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hFCB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFCC} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b001, 12'hFCD} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hFCF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFD0} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b001, 12'hFD1} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hFD3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFD4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b001, 12'hFD5} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hFD6} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b001, 12'hFD7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFD8} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b001, 12'hFD9} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b001, 12'hFDB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b001, 12'hFDC} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b001, 12'hFDD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b001, 12'hFDE} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b001, 12'hFE0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b001, 12'hFE4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b001, 12'hFE8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b001, 12'hFEC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b001, 12'hFF0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b001, 12'hFF4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b001, 12'hFF8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b001, 12'hFFC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b010, 12'h000} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b010, 12'h001} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h003} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h004} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h005} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h008} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h009} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h00A} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h00B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h00D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h00F} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h011} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h012} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h015} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h016} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b010, 12'h017} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b010, 12'h019} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h01C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h01D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h01E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h021} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h025} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h026} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b010, 12'h027} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b010, 12'h029} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h02B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h02D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b010, 12'h02F} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h031} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h033} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h035} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h037} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h038} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b010, 12'h039} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b010, 12'h03B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h03C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h03D} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b010, 12'h03F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h040} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h041} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h043} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h044} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b010, 12'h045} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h047} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h048} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h049} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h04C} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b010, 12'h04D} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h04E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h04F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h050} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h051} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b010, 12'h052} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h059} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h05A} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h05B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h05D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h05F} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h060} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h061} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b010, 12'h062} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h063} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h065} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b010, 12'h066} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h067} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b010, 12'h06B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h06C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h06D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h06E} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h06F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h070} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b010, 12'h071} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h072} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h073} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h074} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h075} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h077} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h078} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b010, 12'h07B} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b010, 12'h07F} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b010, 12'h083} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b010, 12'h085} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b010, 12'h087} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b010, 12'h088} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h089} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h08B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h08C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b010, 12'h08D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h08E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h091} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h092} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h093} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b010, 12'h094} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h096} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h099} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b010, 12'h09D} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h0A1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h0A3} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h0A4} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b010, 12'h0A5} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b010, 12'h0A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0A8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h0A9} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b010, 12'h0AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0AC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h0AD} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h0AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0B0} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b010, 12'h0B4} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b010, 12'h0B8} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b010, 12'h0BD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h0BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0C0} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b010, 12'h0C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h0C2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h0C5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h0C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h0CA} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h0CD} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b010, 12'h0CE} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h0CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0D5} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h0D6} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h0D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0D8} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h0DC} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b010, 12'h0DD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0DE} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h0E0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h0E1} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h0E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0E4} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0E6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0E8} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b010, 12'h0E9} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h0F0} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b010, 12'h0F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h0F2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h0F4} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b010, 12'h0F5} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h0F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0F8} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b010, 12'h0F9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h0FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h0FE} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h100} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b010, 12'h101} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h104} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b010, 12'h105} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h106} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h108} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h109} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h10A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h10D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h10F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h111} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h113} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h115} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h116} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h117} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h11D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h11E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h121} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h122} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h126} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h127} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h12A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h12B} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b010, 12'h132} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h134} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h138} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b010, 12'h139} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h13A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h13C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h13D} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h13F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h141} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h142} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h145} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h148} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h149} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h14A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h14C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h14D} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b010, 12'h14E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h14F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h151} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h153} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h155} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h156} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h159} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h15A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h15B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h15D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h15F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h161} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h162} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h164} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h165} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h166} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h167} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h168} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h16D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h16E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h170} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h171} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h172} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h173} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h174} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'h175} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h176} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h179} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h17A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h17B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h180} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b010, 12'h181} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h182} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h184} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h185} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h188} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h189} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b010, 12'h18C} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b010, 12'h18D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h18E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h190} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h191} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h192} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h193} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h194} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b010, 12'h195} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'h196} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h199} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h19A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h19B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h19C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h19D} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h19F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h1A0} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b010, 12'h1A1} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h1A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h1A4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h1A5} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b010, 12'h1A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h1A8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h1A9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h1AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h1AC} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h1AD} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'h1B6} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h1B8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b010, 12'h1B9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h1BA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h1BD} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b010, 12'h1BE} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h1C1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h1C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h1C6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h1C8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h1C9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h1CA} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h1CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h1CC} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h1CD} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b010, 12'h1CE} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h1CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h1D5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h1D6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h1D8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h1DA} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h1DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h1DC} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b010, 12'h1DD} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'h1E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h1E2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h1E5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h1E6} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h1E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h1E9} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b010, 12'h1EA} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h1ED} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h1F2} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h1F5} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b010, 12'h1F6} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h1F9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h1FC} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b010, 12'h1FD} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h200} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h201} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h203} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h204} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b010, 12'h208} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h209} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h20C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h210} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h211} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h215} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h216} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h218} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b010, 12'h21C} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b010, 12'h220} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b010, 12'h224} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b010, 12'h225} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h226} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h227} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h228} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b010, 12'h22C} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b010, 12'h230} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b010, 12'h234} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b010, 12'h235} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h236} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h237} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h238} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b010, 12'h23C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h23D} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h23E} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h240} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b010, 12'h244} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b010, 12'h246} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h248} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b010, 12'h249} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h24A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h24B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h24C} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'h250} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b010, 12'h254} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b010, 12'h258} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b010, 12'h259} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h25A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h25B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h25C} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'h260} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b010, 12'h264} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b010, 12'h268} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b010, 12'h269} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h26A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h26B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h26C} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b010, 12'h270} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h271} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h272} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h274} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'h278} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b010, 12'h27A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h27C} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b010, 12'h27D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h27E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h27F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h280} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b010, 12'h284} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h285} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h286} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h288} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b010, 12'h28C} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b010, 12'h290} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b010, 12'h291} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h292} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h293} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h294} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b010, 12'h298} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h299} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h29A} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h29C} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b010, 12'h2A0} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b010, 12'h2A4} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b010, 12'h2A5} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h2A6} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h2A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h2A8} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b010, 12'h2AC} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h2AD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h2B0} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b010, 12'h2B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h2B2} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h2B4} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b010, 12'h2B5} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h2B6} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h2B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h2BC} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b010, 12'h2BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h2BE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h2C4} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b010, 12'h2C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h2C6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h2C9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h2CA} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h2D1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h2D2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h2D5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h2D6} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h2DC} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h2DD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h2DE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h2E2} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h2E8} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b010, 12'h2E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h2EA} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h2F0} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b010, 12'h2F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h2F2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h2F4} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b010, 12'h2F5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h2F6} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h2F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h2F8} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b010, 12'h2F9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h2FC} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b010, 12'h2FD} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h300} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h305} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b010, 12'h307} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h309} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h30A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h30D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h30E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h30F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h316} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h319} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b010, 12'h31B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h31C} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b010, 12'h31D} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h31E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h321} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b010, 12'h323} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h324} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b010, 12'h325} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h326} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h329} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b010, 12'h32B} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h32C} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h32D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h32E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h330} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b010, 12'h331} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'h332} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h333} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h335} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b010, 12'h337} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h338} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h339} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h33B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h33C} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b010, 12'h33D} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b010, 12'h33F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h340} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h341} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b010, 12'h342} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h343} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h345} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h346} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h348} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b010, 12'h349} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b010, 12'h34B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h34C} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h34D} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b010, 12'h34E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h34F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h351} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h352} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h354} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b010, 12'h355} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b010, 12'h357} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h358} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b010, 12'h359} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b010, 12'h35A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h35B} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h35C} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h35D} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b010, 12'h35E} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h35F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h361} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h362} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h364} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b010, 12'h365} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h368} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b010, 12'h369} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h36A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h36B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h36C} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b010, 12'h36D} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h36E} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b010, 12'h372} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h373} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h375} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h377} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h378} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h379} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b010, 12'h37A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h37B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h37C} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b010, 12'h37D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h37E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h37F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h380} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b010, 12'h381} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h383} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h384} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b010, 12'h385} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h386} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h387} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h389} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h38A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h390} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h391} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h392} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h393} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h394} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b010, 12'h395} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h396} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h39C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b010, 12'h39D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h39E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h39F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3A0} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b010, 12'h3A1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h3A3} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b010, 12'h3A4} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b010, 12'h3A5} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h3A6} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h3A7} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b010, 12'h3A8} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b010, 12'h3A9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h3AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3AC} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b010, 12'h3AD} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b010, 12'h3AE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h3B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h3B2} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h3B4} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h3B9} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b010, 12'h3BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3BC} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b010, 12'h3BF} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b010, 12'h3C0} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b010, 12'h3C1} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b010, 12'h3C5} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h3C6} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h3C9} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b010, 12'h3CB} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h3CD} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h3CE} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h3D0} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b010, 12'h3D1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h3D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b010, 12'h3D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3D4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h3D8} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b010, 12'h3D9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h3DA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3DD} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h3DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3E0} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h3E1} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b010, 12'h3E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3E4} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h3E5} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'h3E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3E8} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h3E9} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h3EA} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'h3EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3EC} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h3EE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h3F0} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h3F1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3F2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h3F4} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b010, 12'h3F5} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'h3F6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h3F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h3F8} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h3FC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h3FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h3FE} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h400} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b010, 12'h404} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h405} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h407} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h409} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h40A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h40B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h40D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h40E} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b010, 12'h410} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h411} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h412} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h416} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h417} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h418} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h419} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h41A} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'h41C} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h41D} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'h41E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h41F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h421} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h422} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h424} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h425} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h426} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h427} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h428} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h429} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h42A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h42D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h42F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h430} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h431} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h432} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h43A} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b010, 12'h43D} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h43E} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b010, 12'h43F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h440} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h441} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b010, 12'h442} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h444} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b010, 12'h445} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h448} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b010, 12'h449} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b010, 12'h44A} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b010, 12'h44B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h44C} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b010, 12'h44D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h44F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h450} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b010, 12'h451} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b010, 12'h452} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h455} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h456} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h458} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h459} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h45D} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b010, 12'h45F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h461} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h463} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h464} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h465} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h467} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h468} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h469} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b010, 12'h46C} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b010, 12'h46D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h46E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h46F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h471} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h473} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h474} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b010, 12'h475} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h477} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h478} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h479} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'h47D} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h47E} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h47F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h481} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h482} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h484} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b010, 12'h485} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h486} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h488} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'h489} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h48A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h48B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h48D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b010, 12'h48E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h495} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b010, 12'h496} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h49C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h49D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h49E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h4A1} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b010, 12'h4A5} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b010, 12'h4A6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h4A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h4A9} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h4AD} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h4AE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h4AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h4B1} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b010, 12'h4B2} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h4B5} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b010, 12'h4B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h4BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h4BE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h4C1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h4C2} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h4C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h4CA} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h4CD} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h4CE} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'h4D4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h4D6} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h4D8} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b010, 12'h4D9} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b010, 12'h4DA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h4DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h4E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h4E2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h4E6} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h4E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h4EC} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b010, 12'h4EE} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h4F1} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h4F5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h4F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h4F9} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h4FE} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h500} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h501} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h502} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h503} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h505} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h507} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h508} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h50A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h511} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h512} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h515} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h516} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h517} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h51D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h51E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h521} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h522} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h523} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h524} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h525} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h527} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h528} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b010, 12'h529} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b010, 12'h52A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h52B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h52C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h530} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b010, 12'h532} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h535} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h537} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h539} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b010, 12'h53A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h53D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b010, 12'h53E} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'h544} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h546} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h548} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b010, 12'h549} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'h54A} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'h552} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h55A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h560} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h562} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h564} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h565} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h567} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h569} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h56A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h56C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h56D} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h56E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h56F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h570} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'h571} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h572} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h575} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h576} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h577} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h57C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h57D} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b010, 12'h57E} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h580} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b010, 12'h581} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h582} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h584} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h585} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b010, 12'h588} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b010, 12'h589} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h58A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h58D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h58E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h58F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h590} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h594} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h595} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'h597} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h598} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b010, 12'h599} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h59A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h59C} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b010, 12'h59D} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b010, 12'h59E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h59F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h5A6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h5A8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h5A9} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h5AA} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h5AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5AC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b010, 12'h5AD} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'h5AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5B0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h5B1} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h5B2} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h5B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5B4} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b010, 12'h5B5} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5B8} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b010, 12'h5BA} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h5BC} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b010, 12'h5BD} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h5BE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h5BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5C1} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h5C2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5C5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h5C6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5C8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h5CC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h5CD} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'h5CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5D1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h5D2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h5D5} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h5D6} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h5D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5D9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h5DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5DD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h5DE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h5E1} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h5E5} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h5E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5E9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h5EA} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h5EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h5F2} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h5F8} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b010, 12'h5FA} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h5FC} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b010, 12'h601} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h602} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h604} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h605} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b010, 12'h606} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h607} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h608} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h609} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'h60B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h60C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b010, 12'h60D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h610} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b010, 12'h611} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h612} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h613} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h614} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b010, 12'h615} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h616} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h618} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h61D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h61F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h620} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h621} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b010, 12'h622} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h623} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h624} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b010, 12'h625} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h626} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h627} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h629} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h62B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h62C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b010, 12'h62D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h630} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b010, 12'h631} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h632} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h633} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h635} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h636} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h63C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h63D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h63E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h63F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h640} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b010, 12'h641} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h642} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h648} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'h649} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h64A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h64B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h64C} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b010, 12'h64E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h64F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h650} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b010, 12'h652} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b010, 12'h65A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h65D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h65E} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h660} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b010, 12'h662} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h663} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h664} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b010, 12'h666} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b010, 12'h66C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h66D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h66E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h675} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h676} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h679} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h67A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h67B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h67C} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'h67D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h67F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h681} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h683} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h684} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b010, 12'h685} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h686} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b010, 12'h687} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b010, 12'h688} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'h689} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h68B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h68D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h68E} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h691} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h693} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h694} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b010, 12'h695} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h696} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b010, 12'h697} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b010, 12'h698} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'h699} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h69B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h69D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h69F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6A0} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b010, 12'h6A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6A2} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b010, 12'h6A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6A4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h6A6} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h6A8} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'h6A9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h6AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6AE} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h6B1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h6B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6B4} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b010, 12'h6B5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6B6} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b010, 12'h6B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6B8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h6BA} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h6BD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h6BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6C1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h6C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6C4} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h6C6} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h6C8} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b010, 12'h6C9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6CA} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'h6CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6CC} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b010, 12'h6CE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6D2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6D5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6D6} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h6D7} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h6D8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h6DA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6DC} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b010, 12'h6DE} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h6DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6E0} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b010, 12'h6E1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6E2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6E3} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b010, 12'h6E6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6E7} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b010, 12'h6EC} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b010, 12'h6ED} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b010, 12'h6EE} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'h6F0} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'h6F1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h6F3} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b010, 12'h6F4} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b010, 12'h6FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h6FE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h701} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h702} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b010, 12'h703} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h708} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h70A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h711} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h712} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h715} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b010, 12'h716} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b010, 12'h717} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h71C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h71E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h720} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h722} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h724} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b010, 12'h725} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b010, 12'h72A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h72B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h72C} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b010, 12'h72D} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h72E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h730} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'h731} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h732} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h733} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b010, 12'h735} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h739} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h73A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h73E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h73F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h740} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h742} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h744} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b010, 12'h745} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h746} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h74E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h750} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b010, 12'h752} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h753} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h754} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b010, 12'h756} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b010, 12'h75E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h761} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h762} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h76A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h76C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b010, 12'h771} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h773} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h775} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h777} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h779} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h77B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h77D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h77F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h780} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'h782} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h784} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b010, 12'h785} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h786} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h787} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h788} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b010, 12'h789} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b010, 12'h78B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h78C} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b010, 12'h78D} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h78E} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h791} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h792} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h793} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h794} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h796} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h798} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b010, 12'h799} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b010, 12'h79A} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b010, 12'h79B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h79D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h79F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7A1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h7A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7A5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b010, 12'h7A6} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b010, 12'h7A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7A9} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h7AA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b010, 12'h7AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7AE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7B0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b010, 12'h7B1} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b010, 12'h7B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7B4} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b010, 12'h7B5} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h7B6} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h7B9} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h7BA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7BC} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7BE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7C0} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b010, 12'h7C1} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'h7C2} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h7C5} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h7C6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7C8} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'h7CA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7CC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b010, 12'h7CE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h7CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7D0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b010, 12'h7D2} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b010, 12'h7D9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h7DA} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h7DD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h7DE} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h7E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h7E6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h7E9} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h7EA} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h7EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7EC} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b010, 12'h7ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h7EE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7F0} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b010, 12'h7F1} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h7F6} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b010, 12'h7F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'h7F9} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h7FD} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b010, 12'h7FE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'h801} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h802} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h804} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'h80A} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b010, 12'h80E} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b010, 12'h810} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h812} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'h814} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'h818} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b010, 12'h81C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b010, 12'h820} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b010, 12'h824} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'h828} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'h82C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'h830} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'h834} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'h838} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'h83C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'h840} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'h844} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b010, 12'h848} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b010, 12'h84C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b010, 12'h850} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b010, 12'h854} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b010, 12'h858} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b010, 12'h85C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'h860} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b010, 12'h864} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b010, 12'h868} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b010, 12'h86C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b010, 12'h870} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'h874} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'h878} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b010, 12'h87C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b010, 12'h880} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'h884} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b010, 12'h888} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b010, 12'h88C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b010, 12'h890} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b010, 12'h894} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'h898} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b010, 12'h89C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b010, 12'h8A0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b010, 12'h8A4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b010, 12'h8A8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b010, 12'h8AC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b010, 12'h8B0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b010, 12'h8B4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b010, 12'h8B8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b010, 12'h8BC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'h8C0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b010, 12'h8C4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b010, 12'h8C8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b010, 12'h8CC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b010, 12'h8D0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b010, 12'h8D4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b010, 12'h8D8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b010, 12'h8DC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b010, 12'h8E0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b010, 12'h8E4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b010, 12'h8E8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b010, 12'h8EC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b010, 12'h8F0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b010, 12'h8F4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b010, 12'h8F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b010, 12'h8FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b010, 12'h900} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b010, 12'h904} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b010, 12'h908} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b010, 12'h90C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b010, 12'h910} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b010, 12'h914} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b010, 12'h918} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b010, 12'h91C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b010, 12'h920} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b010, 12'h924} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b010, 12'h928} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b010, 12'h92C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b010, 12'h930} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b010, 12'h934} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b010, 12'h938} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b010, 12'h93C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b010, 12'h940} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b010, 12'h944} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b010, 12'h948} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b010, 12'h94C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b010, 12'h950} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b010, 12'h954} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b010, 12'h958} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b010, 12'h95C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b010, 12'h960} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b010, 12'h964} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b010, 12'h968} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b010, 12'h96C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b010, 12'h970} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b010, 12'h974} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b010, 12'h978} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b010, 12'h97C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b010, 12'h980} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'h984} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b010, 12'h988} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b010, 12'h98C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b010, 12'h990} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b010, 12'h994} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'h998} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b010, 12'h99C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b010, 12'h9A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b010, 12'h9A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b010, 12'h9A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b010, 12'h9AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b010, 12'h9B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b010, 12'h9B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b010, 12'h9B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b010, 12'h9BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b010, 12'h9C0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b010, 12'h9C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b010, 12'h9C8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b010, 12'h9CC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b010, 12'h9D0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b010, 12'h9D4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b010, 12'h9D8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b010, 12'h9DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b010, 12'h9E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b010, 12'h9E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b010, 12'h9E8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b010, 12'h9EC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b010, 12'h9F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b010, 12'h9F4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b010, 12'h9F8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b010, 12'h9FC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b010, 12'hA00} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'hA04} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b010, 12'hA08} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b010, 12'hA0C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b010, 12'hA10} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b010, 12'hA14} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hA18} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b010, 12'hA1C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b010, 12'hA20} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b010, 12'hA24} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'hA28} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b010, 12'hA2C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b010, 12'hA30} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b010, 12'hA34} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b010, 12'hA38} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hA3C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'hA40} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b010, 12'hA44} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b010, 12'hA48} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b010, 12'hA4C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b010, 12'hA50} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b010, 12'hA54} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b010, 12'hA58} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b010, 12'hA5C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b010, 12'hA60} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b010, 12'hA64} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b010, 12'hA68} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b010, 12'hA6C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b010, 12'hA70} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b010, 12'hA74} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b010, 12'hA78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b010, 12'hA7C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b010, 12'hA80} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'hA84} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b010, 12'hA88} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b010, 12'hA8C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b010, 12'hA90} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b010, 12'hA94} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b010, 12'hA98} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b010, 12'hA9C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b010, 12'hAA0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b010, 12'hAA4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b010, 12'hAA8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b010, 12'hAAC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b010, 12'hAB0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b010, 12'hAB4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b010, 12'hAB8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b010, 12'hABC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'hAC0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hAC4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b010, 12'hAC8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b010, 12'hACC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b010, 12'hAD0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b010, 12'hAD4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b010, 12'hAD8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b010, 12'hADC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b010, 12'hAE0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b010, 12'hAE4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b010, 12'hAE8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b010, 12'hAEC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b010, 12'hAF0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b010, 12'hAF4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b010, 12'hAF8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b010, 12'hAFC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b010, 12'hB00} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'hB04} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b010, 12'hB08} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b010, 12'hB0C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b010, 12'hB10} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b010, 12'hB14} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b010, 12'hB18} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b010, 12'hB1C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b010, 12'hB20} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b010, 12'hB24} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b010, 12'hB28} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b010, 12'hB2C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b010, 12'hB30} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b010, 12'hB34} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b010, 12'hB38} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b010, 12'hB3C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b010, 12'hB40} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b010, 12'hB44} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b010, 12'hB48} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b010, 12'hB4C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b010, 12'hB50} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b010, 12'hB54} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b010, 12'hB58} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b010, 12'hB5C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b010, 12'hB60} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b010, 12'hB64} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b010, 12'hB68} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b010, 12'hB6C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b010, 12'hB70} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b010, 12'hB74} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b010, 12'hB78} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b010, 12'hB7C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b010, 12'hB80} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b010, 12'hB84} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b010, 12'hB88} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b010, 12'hB8C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b010, 12'hB90} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b010, 12'hB94} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b010, 12'hB98} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b010, 12'hB9C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b010, 12'hBA0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b010, 12'hBA4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b010, 12'hBA8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b010, 12'hBAC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b010, 12'hBB0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b010, 12'hBB4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b010, 12'hBB8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b010, 12'hBBC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b010, 12'hBC0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b010, 12'hBC4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b010, 12'hBC8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b010, 12'hBCC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b010, 12'hBD0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b010, 12'hBD4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b010, 12'hBD8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b010, 12'hBDC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b010, 12'hBE0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b010, 12'hBE4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b010, 12'hBE8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b010, 12'hBEC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b010, 12'hBF0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b010, 12'hBF4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b010, 12'hBF8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b010, 12'hBFC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b010, 12'hC04} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b010, 12'hC08} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b010, 12'hC0C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b010, 12'hC10} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b010, 12'hC14} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b010, 12'hC18} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b010, 12'hC1C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b010, 12'hC20} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b010, 12'hC24} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'hC28} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b010, 12'hC2C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b010, 12'hC30} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'hC34} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b010, 12'hC38} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b010, 12'hC3C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'hC40} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'hC44} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b010, 12'hC48} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b010, 12'hC4C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b010, 12'hC50} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b010, 12'hC54} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b010, 12'hC58} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b010, 12'hC5C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b010, 12'hC60} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b010, 12'hC64} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b010, 12'hC68} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b010, 12'hC6C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b010, 12'hC70} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'hC74} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'hC78} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b010, 12'hC7C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b010, 12'hC80} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hC84} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b010, 12'hC88} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b010, 12'hC8C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b010, 12'hC90} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b010, 12'hC94} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b010, 12'hC98} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b010, 12'hC9C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b010, 12'hCA0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b010, 12'hCA4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b010, 12'hCA8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b010, 12'hCAC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b010, 12'hCB0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b010, 12'hCB4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b010, 12'hCB8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b010, 12'hCBC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hCC0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b010, 12'hCC4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b010, 12'hCC8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b010, 12'hCCC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b010, 12'hCD0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b010, 12'hCD4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b010, 12'hCD8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b010, 12'hCDC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b010, 12'hCE0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b010, 12'hCE4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b010, 12'hCE8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b010, 12'hCEC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b010, 12'hCF0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b010, 12'hCF4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b010, 12'hCF8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b010, 12'hCFC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b010, 12'hD00} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b010, 12'hD04} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b010, 12'hD08} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b010, 12'hD0C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b010, 12'hD10} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b010, 12'hD14} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b010, 12'hD18} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b010, 12'hD1C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b010, 12'hD20} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b010, 12'hD24} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b010, 12'hD28} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b010, 12'hD2C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b010, 12'hD30} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b010, 12'hD34} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b010, 12'hD38} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b010, 12'hD3C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b010, 12'hD40} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b010, 12'hD44} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b010, 12'hD48} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b010, 12'hD4C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b010, 12'hD50} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b010, 12'hD54} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b010, 12'hD58} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b010, 12'hD5C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b010, 12'hD60} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b010, 12'hD64} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b010, 12'hD68} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b010, 12'hD6C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b010, 12'hD70} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b010, 12'hD74} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b010, 12'hD78} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b010, 12'hD7C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b010, 12'hD80} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b010, 12'hD84} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b010, 12'hD88} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b010, 12'hD8C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b010, 12'hD90} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b010, 12'hD94} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'hD98} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b010, 12'hD9C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b010, 12'hDA0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b010, 12'hDA4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b010, 12'hDA8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b010, 12'hDAC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b010, 12'hDB0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b010, 12'hDB4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b010, 12'hDB8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b010, 12'hDBC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b010, 12'hDC0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b010, 12'hDC4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b010, 12'hDC8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b010, 12'hDCC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b010, 12'hDD0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b010, 12'hDD4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b010, 12'hDD8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b010, 12'hDDC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b010, 12'hDE0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b010, 12'hDE4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b010, 12'hDE8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b010, 12'hDEC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b010, 12'hDF0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b010, 12'hDF4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b010, 12'hDF8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b010, 12'hDFC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b010, 12'hE00} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'hE04} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b010, 12'hE08} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b010, 12'hE0C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b010, 12'hE10} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b010, 12'hE14} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hE18} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b010, 12'hE1C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b010, 12'hE20} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b010, 12'hE24} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'hE28} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b010, 12'hE2C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b010, 12'hE30} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b010, 12'hE34} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b010, 12'hE38} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hE3C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b010, 12'hE40} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b010, 12'hE44} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b010, 12'hE48} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b010, 12'hE4C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b010, 12'hE50} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b010, 12'hE54} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b010, 12'hE58} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b010, 12'hE5C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b010, 12'hE60} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b010, 12'hE64} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b010, 12'hE68} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b010, 12'hE6C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b010, 12'hE70} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b010, 12'hE74} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b010, 12'hE78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b010, 12'hE7C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b010, 12'hE80} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'hE84} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b010, 12'hE88} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b010, 12'hE8C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b010, 12'hE90} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b010, 12'hE94} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b010, 12'hE98} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b010, 12'hE9C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b010, 12'hEA0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b010, 12'hEA4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b010, 12'hEA8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b010, 12'hEAC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b010, 12'hEB0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b010, 12'hEB4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b010, 12'hEB8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b010, 12'hEBC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b010, 12'hEC2} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEC6} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEC8} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b010, 12'hECA} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hECC} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b010, 12'hECE} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hED0} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b010, 12'hED2} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hED4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b010, 12'hED6} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hED8} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b010, 12'hEDA} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEDC} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b010, 12'hEDE} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEE0} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b010, 12'hEE2} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEE4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b010, 12'hEE6} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEE8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b010, 12'hEEA} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEEC} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b010, 12'hEEE} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEF0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b010, 12'hEF2} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEF4} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b010, 12'hEF6} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEF8} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b010, 12'hEFA} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hEFC} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b010, 12'hEFE} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b010, 12'hF00} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b010, 12'hF04} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b010, 12'hF05} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b010, 12'hF06} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'hF07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'hF08} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b010, 12'hF09} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b010, 12'hF0A} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF0C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b010, 12'hF0D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF0E} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF10} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b010, 12'hF11} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b010, 12'hF12} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF14} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b010, 12'hF15} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF16} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF18} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b010, 12'hF19} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF1A} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF1C} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b010, 12'hF1D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF1E} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF20} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b010, 12'hF21} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'hF24} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b010, 12'hF25} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'hF28} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b010, 12'hF29} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'hF2C} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b010, 12'hF2D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b010, 12'hF30} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b010, 12'hF31} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hF32} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'hF34} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b010, 12'hF35} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hF36} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'hF38} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b010, 12'hF39} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hF3A} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'hF3C} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b010, 12'hF3D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hF3E} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b010, 12'hF40} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'hF41} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hF42} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'hF44} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'hF46} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'hF48} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b010, 12'hF49} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF4A} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF4C} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b010, 12'hF4D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF4E} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF50} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b010, 12'hF51} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hF52} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'hF54} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b010, 12'hF55} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF56} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF58} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'hF5A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'hF5C} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b010, 12'hF5D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF5E} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF60} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b010, 12'hF61} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hF62} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'hF64} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'hF66} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'hF68} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b010, 12'hF69} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF6A} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF6C} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b010, 12'hF6D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF6E} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF70} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b010, 12'hF71} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hF72} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b010, 12'hF74} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b010, 12'hF75} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF76} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF78} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b010, 12'hF7A} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b010, 12'hF7C} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b010, 12'hF7D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b010, 12'hF7E} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b010, 12'hF80} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b010, 12'hF84} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b010, 12'hF88} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hF8C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b010, 12'hF90} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b010, 12'hF94} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b010, 12'hF98} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b010, 12'hF9C} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b010, 12'hFA0} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b010, 12'hFA4} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFA8} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFAC} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFB0} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFB4} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFB8} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFBC} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFC0} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b010, 12'hFC1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'hFC2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hFC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'hFC4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b010, 12'hFC5} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'hFC8} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b010, 12'hFCC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b010, 12'hFCD} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b010, 12'hFCE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hFCF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'hFD0} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b010, 12'hFD1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b010, 12'hFD2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b010, 12'hFD3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b010, 12'hFD4} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFD8} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFDC} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFE0} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFE4} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFE8} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFEC} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFF0} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFF4} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFF8} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b010, 12'hFFC} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'h000} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h002} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h004} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h006} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h008} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h00A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h00C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h00E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h010} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h012} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h014} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h016} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h018} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h01A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h01C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h01E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h020} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h021} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h022} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h024} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h025} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h026} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h028} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h029} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h02A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h02C} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h02D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h02E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h030} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h031} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h032} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h034} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h035} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h036} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h038} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h039} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h03A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h03C} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h03D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h03E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h040} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h042} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h044} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h046} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h048} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h04A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h04C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h04E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h050} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b011, 12'h051} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h052} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h053} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h054} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b011, 12'h055} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h056} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h057} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h058} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b011, 12'h059} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h05A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h05B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h05C} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b011, 12'h05D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h05E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h05F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h060} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h061} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h062} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h064} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h065} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h066} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h068} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h069} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h06A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h06C} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h06D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h06E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h070} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h071} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h072} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h074} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h075} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h076} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h078} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h079} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h07A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h07C} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h07D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h07E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h080} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h082} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h084} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h086} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h088} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h08A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h08C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h08E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h090} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h092} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h094} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h096} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h098} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h09A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h09C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h09E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h0A0} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h0A1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0A2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0A4} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h0A5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0A6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0A8} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h0A9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0AA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0AC} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h0AD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0AE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0B0} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h0B1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0B2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0B4} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h0B5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0B6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0B8} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h0B9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0BA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0BC} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h0BD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0BE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0C0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h0C2} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h0C4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h0C6} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h0C8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h0CA} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h0CC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h0CE} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h0D0} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b011, 12'h0D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h0D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h0D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h0D4} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b011, 12'h0D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h0D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h0D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h0D8} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b011, 12'h0D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h0DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h0DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h0DC} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b011, 12'h0DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h0DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h0DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h0E0} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h0E1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0E2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0E4} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h0E5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0E6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0E8} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h0E9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0EA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0EC} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h0ED} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0EE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0F0} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h0F1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0F2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0F4} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h0F5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0F6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0F8} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h0F9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0FA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h0FC} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h0FD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h0FE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h100} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h102} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h104} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h106} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h108} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h10A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h10C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h10E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h110} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h112} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h114} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h116} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h118} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h11A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h11C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h11E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h120} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h121} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h122} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h124} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h125} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h126} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h128} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h129} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h12A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h12C} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h12D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h12E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h130} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h131} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h132} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h134} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h135} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h136} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h138} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h139} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h13A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h13C} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h13D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h13E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h140} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h142} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h144} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h146} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h148} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h14A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h14C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h14E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h150} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b011, 12'h151} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h152} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h153} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h154} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b011, 12'h155} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h156} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h157} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h158} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b011, 12'h159} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h15A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h15B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h15C} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b011, 12'h15D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h15E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h15F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h160} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h161} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h162} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h164} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h165} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h166} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h168} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h169} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h16A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h16C} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h16D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h16E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h170} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h171} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h172} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h174} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h175} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h176} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h178} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h179} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h17A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h17C} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h17D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h17E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h180} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h182} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h184} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h186} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h188} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h18A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h18C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h18E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h190} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h192} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h194} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h196} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h198} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h19A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h19C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h19E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h1A0} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h1A1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1A2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1A4} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h1A5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1A6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1A8} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h1A9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1AA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1AC} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h1AD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1AE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1B0} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h1B1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1B2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1B4} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h1B5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1B6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1B8} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h1B9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1BA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1BC} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'h1BD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1BE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1C0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h1C2} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h1C4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h1C6} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h1C8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h1CA} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h1CC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'h1CE} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h1D0} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b011, 12'h1D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h1D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h1D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h1D4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b011, 12'h1D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h1D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h1D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h1D8} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b011, 12'h1D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h1DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h1DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h1DC} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b011, 12'h1DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h1DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h1DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h1E0} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h1E1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1E2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1E4} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h1E5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1E6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1E8} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h1E9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1EA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1EC} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h1ED} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1EE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1F0} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h1F1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1F2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1F4} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h1F5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1F6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1F8} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h1F9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1FA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h1FC} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b011, 12'h1FD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h1FE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h200} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h202} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h204} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h206} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h208} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h20A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h20C} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h20E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h210} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h212} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h214} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h216} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h218} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h21A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h21C} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h21E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h220} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b011, 12'h221} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h222} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h224} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b011, 12'h225} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h226} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h228} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b011, 12'h229} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h22A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h22C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b011, 12'h22D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h22E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h230} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b011, 12'h231} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h232} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h234} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b011, 12'h235} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h236} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h238} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b011, 12'h239} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h23A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h23C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b011, 12'h23D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h23E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h240} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h242} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h244} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h246} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h248} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h24A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h24C} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b011, 12'h24E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h250} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b011, 12'h251} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h252} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h253} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h254} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b011, 12'h255} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h256} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h257} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h258} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b011, 12'h259} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h25A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h25B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h25C} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b011, 12'h25D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h25E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h25F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h260} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b011, 12'h261} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h262} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h264} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b011, 12'h265} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h266} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h268} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b011, 12'h269} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h26A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h26C} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b011, 12'h26D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h26E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h270} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b011, 12'h271} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h272} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h274} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b011, 12'h275} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h276} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h278} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b011, 12'h279} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h27A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h27C} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b011, 12'h27D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h27E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h280} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h281} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h282} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h284} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h285} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h286} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h288} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h289} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h28A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h28C} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h28D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h28E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h290} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h291} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h292} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h294} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h295} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h296} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h298} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h299} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h29A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h29C} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h29D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h29E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h2A0} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b011, 12'h2A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2A2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2A4} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b011, 12'h2A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2A6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2A8} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b011, 12'h2A9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2AA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2AC} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b011, 12'h2AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2AE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2B0} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b011, 12'h2B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2B2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2B4} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b011, 12'h2B5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2B6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2B8} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b011, 12'h2B9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2BA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2BC} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b011, 12'h2BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2BE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2C0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h2C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2C2} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h2C4} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h2C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2C6} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h2C8} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h2C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2CA} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h2CC} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b011, 12'h2CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2CE} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h2D0} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b011, 12'h2D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h2D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h2D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h2D4} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b011, 12'h2D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h2D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h2D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h2D8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b011, 12'h2D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h2DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h2DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h2DC} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b011, 12'h2DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h2DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h2DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h2E0} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b011, 12'h2E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2E2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2E4} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b011, 12'h2E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2E6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2E8} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b011, 12'h2E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2EA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2EC} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b011, 12'h2ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2EE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2F0} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b011, 12'h2F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2F2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2F4} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b011, 12'h2F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2F6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2F8} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b011, 12'h2F9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2FA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h2FC} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b011, 12'h2FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h2FE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h300} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h302} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h304} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h306} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h308} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h30A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h30C} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h30E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h310} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h312} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h314} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h316} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h318} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h31A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h31C} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h31E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h320} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b011, 12'h321} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h322} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h324} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b011, 12'h325} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h326} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h328} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b011, 12'h329} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h32A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h32C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b011, 12'h32D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h32E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h330} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b011, 12'h331} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h332} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h334} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b011, 12'h335} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h336} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h338} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b011, 12'h339} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h33A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h33C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b011, 12'h33D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h33E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h340} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h342} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h344} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h346} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h348} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h34A} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h34C} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b011, 12'h34E} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b011, 12'h350} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b011, 12'h351} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h352} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h353} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h354} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b011, 12'h355} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h356} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h357} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h358} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b011, 12'h359} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h35A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h35B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h35C} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b011, 12'h35D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h35E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h35F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h360} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b011, 12'h361} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h362} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h364} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b011, 12'h365} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h366} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h368} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b011, 12'h369} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h36A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h36C} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b011, 12'h36D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h36E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h370} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b011, 12'h371} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h372} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h374} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b011, 12'h375} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h376} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h378} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b011, 12'h379} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h37A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h37C} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b011, 12'h37D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b011, 12'h37E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h380} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h381} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h382} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h384} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h385} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h386} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h388} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h389} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h38A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h38C} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h38D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h38E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h390} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h391} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h392} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h394} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h395} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h396} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h398} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h399} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h39A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h39C} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h39D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h39E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h3A0} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b011, 12'h3A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3A2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3A4} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b011, 12'h3A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3A6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3A8} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b011, 12'h3A9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3AA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3AC} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b011, 12'h3AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3AE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3B0} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b011, 12'h3B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3B2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3B4} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b011, 12'h3B5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3B6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3B8} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b011, 12'h3B9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3BA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3BC} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b011, 12'h3BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3BE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3C0} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h3C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3C2} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h3C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h3C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3C6} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h3C8} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h3C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3CA} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h3CC} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b011, 12'h3CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3CE} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h3D0} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b011, 12'h3D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h3D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h3D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h3D4} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b011, 12'h3D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h3D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h3D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h3D8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b011, 12'h3D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h3DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h3DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h3DC} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b011, 12'h3DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h3DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h3DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h3E0} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b011, 12'h3E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3E2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3E4} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b011, 12'h3E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3E6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3E8} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b011, 12'h3E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3EA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3EC} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b011, 12'h3ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3EE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3F0} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b011, 12'h3F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3F2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3F4} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b011, 12'h3F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3F6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3F8} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b011, 12'h3F9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3FA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h3FC} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b011, 12'h3FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h3FE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h400} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h401} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h402} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h404} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h405} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h406} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h408} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h409} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h40A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h40C} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h40D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h40E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h410} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h411} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h412} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h414} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h415} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h416} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h418} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h419} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h41A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h41C} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h41D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h41E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h420} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b011, 12'h421} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h422} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h424} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b011, 12'h425} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h426} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h428} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b011, 12'h429} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h42A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h42C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b011, 12'h42D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h42E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h430} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b011, 12'h431} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h432} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h434} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b011, 12'h435} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h436} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h438} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b011, 12'h439} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h43A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h43C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b011, 12'h43D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h43E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h440} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h441} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h442} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h444} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h445} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h446} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h448} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h449} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h44A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h44C} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b011, 12'h44D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h44E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h450} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b011, 12'h451} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h452} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h453} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h454} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b011, 12'h455} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h456} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h457} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h458} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b011, 12'h459} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h45A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h45B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h45C} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b011, 12'h45D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h45E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h45F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h460} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b011, 12'h461} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h462} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h464} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b011, 12'h465} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h466} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h468} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b011, 12'h469} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h46A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h46C} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b011, 12'h46D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h46E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h470} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b011, 12'h471} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h472} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h474} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b011, 12'h475} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h476} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h478} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b011, 12'h479} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h47A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h47C} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b011, 12'h47D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h47E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h480} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h481} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h482} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h484} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h485} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h486} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h488} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h489} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h48A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h48C} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h48D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h48E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h490} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h491} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h492} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h494} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h495} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h496} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h498} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h499} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h49A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h49C} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h49D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h49E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h4A0} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b011, 12'h4A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4A2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4A4} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b011, 12'h4A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4A6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4A8} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b011, 12'h4A9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4AA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4AC} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b011, 12'h4AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4AE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4B0} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b011, 12'h4B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4B2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4B4} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b011, 12'h4B5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4B6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4B8} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b011, 12'h4B9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4BA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4BC} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b011, 12'h4BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4BE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4C0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h4C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4C2} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h4C4} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h4C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4C6} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h4C8} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h4C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4CA} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h4CC} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b011, 12'h4CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4CE} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h4D0} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b011, 12'h4D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h4D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h4D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h4D4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b011, 12'h4D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h4D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h4D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h4D8} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b011, 12'h4D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h4DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h4DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h4DC} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b011, 12'h4DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h4DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h4DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h4E0} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b011, 12'h4E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4E2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4E4} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b011, 12'h4E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4E6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4E8} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b011, 12'h4E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4EA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4EC} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b011, 12'h4ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4EE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4F0} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b011, 12'h4F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4F2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4F4} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b011, 12'h4F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4F6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4F8} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b011, 12'h4F9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4FA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h4FC} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b011, 12'h4FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h4FE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h500} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h501} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h502} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h504} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h505} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h506} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h508} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h509} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h50A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h50C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h50D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h50E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h510} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h511} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h512} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h514} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h515} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h516} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h518} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h519} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h51A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h51C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h51D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h51E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h520} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b011, 12'h521} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h522} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h524} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b011, 12'h525} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h526} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h528} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b011, 12'h529} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h52A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h52C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b011, 12'h52D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h52E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h530} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b011, 12'h531} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h532} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h534} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b011, 12'h535} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h536} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h538} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b011, 12'h539} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h53A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h53C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b011, 12'h53D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h53E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h540} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h541} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h542} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h544} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h545} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h546} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h548} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h549} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h54A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h54C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h54D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h54E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h550} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b011, 12'h551} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h552} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h553} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h554} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b011, 12'h555} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h556} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h557} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h558} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b011, 12'h559} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h55A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h55B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h55C} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b011, 12'h55D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h55E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h55F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h560} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b011, 12'h561} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h562} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h564} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b011, 12'h565} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h566} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h568} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b011, 12'h569} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h56A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h56C} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b011, 12'h56D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h56E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h570} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b011, 12'h571} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h572} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h574} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b011, 12'h575} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h576} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h578} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b011, 12'h579} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h57A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h57C} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b011, 12'h57D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h57E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h580} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h581} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h582} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h584} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h585} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h586} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h588} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h589} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h58A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h58C} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h58D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h58E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h590} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h591} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h592} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h594} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h595} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h596} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h598} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h599} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h59A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h59C} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h59D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h59E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h5A0} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b011, 12'h5A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5A2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5A4} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b011, 12'h5A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5A6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5A8} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b011, 12'h5A9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5AA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5AC} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b011, 12'h5AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5AE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5B0} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b011, 12'h5B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5B2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5B4} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b011, 12'h5B5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5B6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5B8} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b011, 12'h5B9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5BA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5BC} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b011, 12'h5BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5BE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5C0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h5C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5C2} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h5C4} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h5C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5C6} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h5C8} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h5C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5CA} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h5CC} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b011, 12'h5CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5CE} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h5D0} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b011, 12'h5D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h5D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h5D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h5D4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b011, 12'h5D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h5D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h5D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h5D8} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b011, 12'h5D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h5DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h5DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h5DC} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b011, 12'h5DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h5DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h5DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h5E0} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b011, 12'h5E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5E2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5E4} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b011, 12'h5E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5E6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5E8} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b011, 12'h5E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5EA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5EC} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b011, 12'h5ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5EE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5F0} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b011, 12'h5F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5F2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5F4} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b011, 12'h5F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5F6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5F8} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b011, 12'h5F9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5FA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h5FC} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b011, 12'h5FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h5FE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h600} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h601} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h602} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h604} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h605} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h606} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h608} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h609} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h60A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h60C} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h60D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h60E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h610} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h611} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h612} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h614} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h615} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h616} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h618} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h619} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h61A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h61C} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h61D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h61E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h620} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'h621} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h622} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h624} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'h625} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h626} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h628} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'h629} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h62A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h62C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'h62D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h62E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h630} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'h631} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h632} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h634} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'h635} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h636} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h638} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'h639} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h63A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h63C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'h63D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h63E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h640} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h641} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h642} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h644} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h645} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h646} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h648} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h649} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h64A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h64C} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b011, 12'h64D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h64E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h650} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b011, 12'h651} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h652} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h653} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h654} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b011, 12'h655} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h656} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h657} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h658} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b011, 12'h659} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h65A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h65B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h65C} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b011, 12'h65D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h65E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h65F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h660} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b011, 12'h661} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h662} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h664} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b011, 12'h665} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h666} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h668} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b011, 12'h669} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h66A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h66C} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b011, 12'h66D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h66E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h670} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b011, 12'h671} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h672} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h674} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b011, 12'h675} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h676} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h678} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b011, 12'h679} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h67A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h67C} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b011, 12'h67D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h67E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h680} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h681} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h682} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h684} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h685} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h686} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h688} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h689} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h68A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h68C} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h68D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h68E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h690} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h691} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h692} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h694} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h695} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h696} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h698} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h699} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h69A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h69C} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h69D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h69E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h6A0} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b011, 12'h6A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6A2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6A4} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b011, 12'h6A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6A6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6A8} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b011, 12'h6A9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6AA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6AC} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b011, 12'h6AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6AE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6B0} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b011, 12'h6B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6B2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6B4} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b011, 12'h6B5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6B6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6B8} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b011, 12'h6B9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6BA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6BC} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b011, 12'h6BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6BE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6C0} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h6C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6C2} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h6C4} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h6C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6C6} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h6C8} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h6C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6CA} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h6CC} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h6CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6CE} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h6D0} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b011, 12'h6D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h6D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h6D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h6D4} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b011, 12'h6D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h6D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h6D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h6D8} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b011, 12'h6D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h6DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h6DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h6DC} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b011, 12'h6DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h6DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h6DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h6E0} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b011, 12'h6E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6E2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6E4} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b011, 12'h6E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6E6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6E8} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b011, 12'h6E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6EA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6EC} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b011, 12'h6ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6EE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6F0} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b011, 12'h6F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6F2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6F4} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b011, 12'h6F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6F6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6F8} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b011, 12'h6F9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6FA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h6FC} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b011, 12'h6FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h6FE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h700} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h701} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h702} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h704} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h705} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h706} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h708} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h709} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h70A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h70C} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h70D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h70E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h710} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h711} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h712} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h714} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h715} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h716} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h718} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h719} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h71A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h71C} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h71D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h71E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h720} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'h721} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h722} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h724} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'h725} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h726} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h728} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'h729} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h72A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h72C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'h72D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h72E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h730} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'h731} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h732} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h734} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'h735} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h736} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h738} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'h739} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h73A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h73C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'h73D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h73E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h740} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h741} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h742} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h744} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h745} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h746} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h748} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h749} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h74A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h74C} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b011, 12'h74D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h74E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h750} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b011, 12'h751} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h752} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h753} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h754} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b011, 12'h755} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h756} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h757} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h758} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b011, 12'h759} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h75A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h75B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h75C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b011, 12'h75D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h75E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h75F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h760} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b011, 12'h761} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h762} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h764} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b011, 12'h765} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h766} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h768} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b011, 12'h769} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h76A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h76C} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b011, 12'h76D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h76E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h770} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b011, 12'h771} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h772} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h774} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b011, 12'h775} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h776} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h778} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b011, 12'h779} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h77A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h77C} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b011, 12'h77D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h77E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h780} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h781} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h782} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h784} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h785} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h786} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h788} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h789} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h78A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h78C} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h78D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h78E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h790} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h791} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h792} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h794} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h795} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h796} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h798} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h799} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h79A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h79C} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h79D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h79E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h7A0} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b011, 12'h7A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7A2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7A4} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b011, 12'h7A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7A6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7A8} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b011, 12'h7A9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7AA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7AC} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b011, 12'h7AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7AE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7B0} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b011, 12'h7B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7B2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7B4} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b011, 12'h7B5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7B6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7B8} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b011, 12'h7B9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7BA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7BC} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b011, 12'h7BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7BE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7C0} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h7C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7C2} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h7C4} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h7C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7C6} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h7C8} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h7C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7CA} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h7CC} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b011, 12'h7CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7CE} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h7D0} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b011, 12'h7D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h7D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h7D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h7D4} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b011, 12'h7D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h7D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h7D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h7D8} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b011, 12'h7D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h7DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h7DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h7DC} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b011, 12'h7DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h7DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h7DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h7E0} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b011, 12'h7E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7E2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7E4} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b011, 12'h7E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7E6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7E8} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b011, 12'h7E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7EA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7EC} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b011, 12'h7ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7EE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7F0} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b011, 12'h7F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7F2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7F4} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b011, 12'h7F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7F6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7F8} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b011, 12'h7F9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7FA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h7FC} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b011, 12'h7FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h7FE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h800} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h801} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h802} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h804} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h805} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h806} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h808} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h809} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h80A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h80C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h80D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h80E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h810} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h811} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h812} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h814} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h815} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h816} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h818} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h819} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h81A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h81C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h81D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h81E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h820} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h821} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h822} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h824} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h825} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h826} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h828} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h829} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h82A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h82C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h82D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h82E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h830} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h831} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h832} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h834} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h835} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h836} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h838} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h839} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h83A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h83C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h83D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h83E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h840} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h841} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h842} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h844} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h845} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h846} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h848} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h849} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h84A} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h84C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h84D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h84E} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'h850} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b011, 12'h851} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h852} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h853} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h854} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b011, 12'h855} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h856} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h857} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h858} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b011, 12'h859} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h85A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h85B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h85C} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b011, 12'h85D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h85E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h85F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h860} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h861} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h862} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h864} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h865} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h866} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h868} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h869} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h86A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h86C} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h86D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h86E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h870} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h871} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h872} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h874} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h875} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h876} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h878} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h879} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h87A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h87C} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h87D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h87E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'h880} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h881} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h882} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h883} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h884} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h885} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h886} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h887} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h888} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h889} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h88A} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h88B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h88C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h88D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h88E} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h88F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h890} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h891} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h892} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h893} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h894} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h895} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h896} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h897} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h898} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h899} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h89A} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h89B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h89C} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h89D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h89E} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h89F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8A0} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h8A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8A2} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8A4} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h8A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8A6} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8A8} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h8A9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8AA} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8AC} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h8AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8AE} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8B0} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h8B1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8B2} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8B4} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h8B5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8B6} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8B8} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h8B9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8BA} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8BC} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b011, 12'h8BD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8BE} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8C0} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h8C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8C2} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h8C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8C4} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h8C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8C6} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h8C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8C8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h8C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8CA} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h8CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8CC} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b011, 12'h8CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8CE} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h8CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8D0} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b011, 12'h8D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h8D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h8D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8D4} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b011, 12'h8D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h8D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h8D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8D8} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b011, 12'h8D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h8DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h8DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8DC} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b011, 12'h8DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h8DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h8DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8E0} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h8E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8E2} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8E4} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h8E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8E6} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8E8} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h8E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8EA} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8EC} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h8ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8EE} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8F0} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h8F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8F2} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8F4} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h8F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8F6} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8F8} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h8F9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8FA} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h8FC} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b011, 12'h8FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'h8FE} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h8FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h900} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h901} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h902} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h903} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h904} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h905} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h906} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h907} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h908} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h909} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h90A} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h90B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h90C} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h90D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h90E} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h90F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h910} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h911} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h912} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h913} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h914} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h915} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h916} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h917} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h918} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h919} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h91A} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h91B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h91C} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h91D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h91E} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h91F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h920} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b011, 12'h921} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h922} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h923} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h924} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b011, 12'h925} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h926} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h927} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h928} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b011, 12'h929} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h92A} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h92B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h92C} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b011, 12'h92D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h92E} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h92F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h930} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b011, 12'h931} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h932} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h933} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h934} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b011, 12'h935} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h936} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h937} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h938} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b011, 12'h939} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h93A} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h93B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h93C} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b011, 12'h93D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h93E} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h93F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h940} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h941} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h942} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h943} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h944} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h945} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h946} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h947} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h948} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h949} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h94A} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h94B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h94C} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'h94D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h94E} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h94F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h950} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b011, 12'h951} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h952} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h953} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h954} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b011, 12'h955} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h956} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h957} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h958} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b011, 12'h959} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h95A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h95B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h95C} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b011, 12'h95D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h95E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h95F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h960} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b011, 12'h961} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h962} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h963} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h964} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b011, 12'h965} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h966} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h967} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h968} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b011, 12'h969} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h96A} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h96B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h96C} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b011, 12'h96D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h96E} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h96F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h970} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b011, 12'h971} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h972} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h973} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h974} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b011, 12'h975} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h976} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h977} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h978} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b011, 12'h979} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h97A} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h97B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h97C} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b011, 12'h97D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h97E} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h97F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h980} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h981} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h982} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h983} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h984} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h985} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h986} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h987} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h988} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h989} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h98A} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h98B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h98C} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h98D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h98E} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h98F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h990} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h991} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h992} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h993} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h994} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h995} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h996} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h997} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h998} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h999} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h99A} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h99B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h99C} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h99D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h99E} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h99F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9A0} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b011, 12'h9A1} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9A2} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9A4} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b011, 12'h9A5} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9A6} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9A8} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b011, 12'h9A9} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9AA} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9AC} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b011, 12'h9AD} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9AE} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9B0} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b011, 12'h9B1} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9B2} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9B4} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b011, 12'h9B5} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9B6} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9B8} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b011, 12'h9B9} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9BA} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9BC} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b011, 12'h9BD} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9BE} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9C0} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h9C1} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9C2} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h9C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9C4} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h9C5} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9C6} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h9C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9C8} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h9C9} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9CA} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h9CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9CC} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b011, 12'h9CD} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9CE} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'h9CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9D0} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b011, 12'h9D1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h9D2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h9D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9D4} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b011, 12'h9D5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h9D6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h9D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9D8} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b011, 12'h9D9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h9DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h9DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9DC} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b011, 12'h9DD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'h9DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'h9DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9E0} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b011, 12'h9E1} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9E2} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9E4} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b011, 12'h9E5} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9E6} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9E8} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b011, 12'h9E9} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9EA} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9EC} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b011, 12'h9ED} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9EE} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9F0} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b011, 12'h9F1} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9F2} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9F4} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b011, 12'h9F5} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9F6} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9F8} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b011, 12'h9F9} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9FA} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'h9FC} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b011, 12'h9FD} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b011, 12'h9FE} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b011, 12'h9FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA00} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA01} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA02} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA04} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA05} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA06} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA08} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA09} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA0A} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA0B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA0C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA0D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA0E} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA0F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA10} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA11} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA12} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA14} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA15} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA16} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA17} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA18} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA19} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA1A} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA1B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA1C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA1D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA1E} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA1F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA20} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b011, 12'hA21} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA22} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA24} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b011, 12'hA25} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA26} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA28} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b011, 12'hA29} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA2A} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA2C} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b011, 12'hA2D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA2E} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA30} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b011, 12'hA31} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA32} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA33} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA34} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b011, 12'hA35} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA36} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA38} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b011, 12'hA39} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA3A} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA3C} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b011, 12'hA3D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA3E} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA40} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA41} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA42} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA44} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA45} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA46} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA47} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA48} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA49} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA4A} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA4C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hA4D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA4E} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b011, 12'hA4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA50} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b011, 12'hA51} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hA52} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hA53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA54} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b011, 12'hA55} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hA56} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hA57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA58} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b011, 12'hA59} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hA5A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hA5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA5C} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b011, 12'hA5D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hA5E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hA5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA60} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b011, 12'hA61} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA62} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA63} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA64} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b011, 12'hA65} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA66} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA68} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b011, 12'hA69} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA6A} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA6C} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b011, 12'hA6D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA6E} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA70} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b011, 12'hA71} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA72} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA74} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b011, 12'hA75} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA76} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA77} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA78} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b011, 12'hA79} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA7A} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA7C} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b011, 12'hA7D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA7E} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b011, 12'hA7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hA81} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA82} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hA85} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA86} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hA89} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA8A} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hA8D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA8E} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hA91} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA92} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hA95} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA96} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hA99} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA9A} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hA9D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hA9E} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hAA0} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hAA1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAA2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAA4} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hAA5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAA6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAA8} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hAA9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAAA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAAC} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hAAD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAAE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAB0} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hAB1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAB2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAB4} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hAB5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAB6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAB8} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hAB9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hABA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hABC} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hABD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hABE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAC1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAC2} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hAC5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAC6} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hAC9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hACA} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hACD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hACE} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hAD0} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b011, 12'hAD1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hAD2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hAD3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hAD4} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b011, 12'hAD5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hAD6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hAD7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hAD8} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b011, 12'hAD9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hADA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hADB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hADC} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b011, 12'hADD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hADE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hADF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hAE0} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hAE1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAE2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAE4} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hAE5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAE6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAE8} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hAE9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAEA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAEC} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hAED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAEE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAF0} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hAF1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAF2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAF4} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hAF5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAF6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAF8} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hAF9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAFA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hAFC} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hAFD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hAFE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hB00} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB01} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB02} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB04} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB05} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB06} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB08} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB09} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB0A} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB0C} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB0D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB0E} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB10} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB11} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB12} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB14} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB15} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB16} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB18} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB19} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB1A} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB1C} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB1D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB1E} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB20} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB21} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB22} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB24} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB25} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB26} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB28} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB29} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB2A} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB2C} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB2D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB2E} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB30} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB31} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB32} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB34} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB35} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB36} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB38} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB39} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB3A} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB3C} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB3D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB3E} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB40} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB41} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hB42} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hB44} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB45} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hB46} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB47} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hB48} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB49} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hB4A} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hB4C} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB4D} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hB4E} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hB50} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB51} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hB52} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hB54} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB55} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hB56} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hB58} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB59} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hB5A} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hB5C} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB5D} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hB5E} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hB60} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB61} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB62} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB64} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB65} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB66} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB68} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB69} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB6A} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB6C} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB6D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB6E} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB70} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB71} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB72} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB74} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB75} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB76} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB78} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB79} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB7A} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB7C} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b011, 12'hB7D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hB7E} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hB81} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hB82} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hB85} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hB86} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hB89} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hB8A} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hB8D} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hB8E} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hB91} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hB92} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hB95} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hB96} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hB99} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hB9A} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hB9D} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hB9E} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hBA0} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hBA1} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBA2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBA4} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hBA5} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBA6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBA8} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hBA9} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBAA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBAC} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hBAD} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBAE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBB0} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hBB1} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBB2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBB4} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hBB5} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBB6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBB8} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hBB9} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBBA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBBC} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b011, 12'hBBD} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBBE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBC1} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBC2} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hBC5} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBC6} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hBC9} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBCA} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hBCD} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBCE} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hBD0} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b011, 12'hBD1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hBD2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hBD3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hBD4} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b011, 12'hBD5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hBD6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hBD7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hBD8} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b011, 12'hBD9} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hBDA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hBDB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hBDC} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b011, 12'hBDD} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b011, 12'hBDE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b011, 12'hBDF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hBE0} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hBE1} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBE2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBE4} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hBE5} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBE6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBE8} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hBE9} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBEA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBEC} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hBED} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBEE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBF0} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hBF1} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBF2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBF4} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hBF5} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBF6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBF8} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hBF9} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBFA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hBFC} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b011, 12'hBFD} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b011, 12'hBFE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hC00} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b011, 12'hC01} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC02} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b011, 12'hC03} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC04} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b011, 12'hC05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hC06} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hC07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hC08} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hC0C} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b011, 12'hC10} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b011, 12'hC11} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC12} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b011, 12'hC13} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC14} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b011, 12'hC18} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b011, 12'hC1C} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b011, 12'hC20} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b011, 12'hC21} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC22} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b011, 12'hC23} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC24} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hC28} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b011, 12'hC2C} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hC30} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b011, 12'hC31} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC32} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b011, 12'hC33} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC34} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hC38} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b011, 12'hC3C} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hC40} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b011, 12'hC41} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC42} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b011, 12'hC43} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC44} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b011, 12'hC45} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC46} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b011, 12'hC47} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b011, 12'hC48} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b011, 12'hC4C} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hC50} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b011, 12'hC51} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC52} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b011, 12'hC53} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC54} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hC58} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b011, 12'hC59} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b011, 12'hC5D} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b011, 12'hC5E} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b011, 12'hC5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hC60} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b011, 12'hC61} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC62} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b011, 12'hC63} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC64} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b011, 12'hC66} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hC68} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b011, 12'hC69} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hC6A} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b011, 12'hC6C} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b011, 12'hC6D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC6E} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b011, 12'hC70} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b011, 12'hC71} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC72} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b011, 12'hC73} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC74} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hC78} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b011, 12'hC79} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b011, 12'hC7A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hC7C} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hC80} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b011, 12'hC83} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b011, 12'hC84} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b011, 12'hC88} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b011, 12'hC8B} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b011, 12'hC8C} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b011, 12'hC90} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hC91} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC92} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hC93} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC94} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hC95} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC96} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hC97} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b011, 12'hC98} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hC99} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC9A} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hC9B} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hC9C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hC9D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hC9E} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hC9F} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b011, 12'hCA0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCA1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCA2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCA3} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hCA4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCA5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCA6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCA7} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b011, 12'hCA8} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hCA9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b011, 12'hCAB} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b011, 12'hCAC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCAD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCAE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCAF} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b011, 12'hCB0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCB1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCB2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCB3} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hCB4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCB5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCB6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCB7} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b011, 12'hCB8} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b011, 12'hCB9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b011, 12'hCBB} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b011, 12'hCBC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCBD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCBE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCBF} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b011, 12'hCC0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCC1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCC2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCC3} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b011, 12'hCC4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCC5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCC6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCC7} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b011, 12'hCC8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCC9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCCA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCCB} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b011, 12'hCCC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCCD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCCE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCCF} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b011, 12'hCD0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCD1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCD2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCD3} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b011, 12'hCD4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCD5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCD6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCD7} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b011, 12'hCD8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCD9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCDA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCDB} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b011, 12'hCDC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCDD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCDE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCDF} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b011, 12'hCE0} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCE1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCE2} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCE3} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b011, 12'hCE4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCE5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCE6} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCE7} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b011, 12'hCE8} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCE9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCEA} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCEB} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b011, 12'hCEC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b011, 12'hCED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCEE} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b011, 12'hCEF} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b011, 12'hCF1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCF2} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b011, 12'hCF5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCF6} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b011, 12'hCF9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCFA} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b011, 12'hCFD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hCFE} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b011, 12'hD00} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b011, 12'hD04} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b011, 12'hD08} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b011, 12'hD0C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b011, 12'hD10} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b011, 12'hD14} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hD18} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hD1C} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b011, 12'hD20} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b011, 12'hD24} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b011, 12'hD28} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b011, 12'hD2C} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b011, 12'hD30} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'hD34} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'hD38} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'hD3C} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b011, 12'hD40} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'hD41} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b011, 12'hD42} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hD43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hD44} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'hD45} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b011, 12'hD46} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hD47} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hD48} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'hD49} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b011, 12'hD4A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hD4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hD4C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b011, 12'hD4D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b011, 12'hD4E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b011, 12'hD4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hD50} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b011, 12'hD54} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b011, 12'hD58} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b011, 12'hD5C} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b011, 12'hD60} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b011, 12'hD62} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b011, 12'hD64} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b011, 12'hD66} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b011, 12'hD68} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b011, 12'hD6A} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b011, 12'hD6C} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b011, 12'hD6E} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b011, 12'hD70} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b011, 12'hD74} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b011, 12'hD78} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b011, 12'hD7C} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b011, 12'hD80} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b011, 12'hD84} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b011, 12'hD88} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b011, 12'hD8C} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b011, 12'hD90} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hD94} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hD98} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b011, 12'hD9C} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b011, 12'hDA0} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b011, 12'hDA4} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b011, 12'hDA8} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b011, 12'hDAC} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b011, 12'hDB0} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hDB4} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hDB8} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b011, 12'hDBC} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b011, 12'hDC0} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b011, 12'hDC4} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b011, 12'hDC8} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b011, 12'hDCC} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b011, 12'hDD0} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hDD4} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hDD8} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b011, 12'hDDC} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b011, 12'hDE0} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b011, 12'hDE4} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b011, 12'hDE8} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b011, 12'hDEC} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b011, 12'hDF0} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hDF4} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b011, 12'hDF8} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b011, 12'hDFC} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b011, 12'hE00} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE04} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE08} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE0C} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE10} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE14} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE18} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE1C} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE20} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE24} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE28} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE2C} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE30} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE34} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE38} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE3C} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE40} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE44} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE48} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE4C} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE50} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE54} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE58} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE5C} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE60} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE64} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE68} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE6C} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE70} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE74} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE78} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE7C} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b011, 12'hE80} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hE84} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hE88} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hE8C} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hE90} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hE94} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hE98} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hE9C} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEA0} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEA4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEA8} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEAC} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEB0} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEB4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEB8} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEBC} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEC0} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEC4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEC8} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hECC} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hED0} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hED4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hED8} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEDC} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEE0} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEE4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEE8} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEEC} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEF0} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEF4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEF8} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hEFC} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b011, 12'hF01} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b011, 12'hF02} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF05} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b011, 12'hF06} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF09} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b011, 12'hF0A} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF0B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF0D} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b011, 12'hF0E} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF0F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF11} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b011, 12'hF12} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF15} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b011, 12'hF16} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF17} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF19} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b011, 12'hF1A} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF1B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF1D} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b011, 12'hF1E} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF1F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF21} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b011, 12'hF22} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF25} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b011, 12'hF26} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF29} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b011, 12'hF2A} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF2D} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b011, 12'hF2E} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF31} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hF32} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF33} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF35} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hF36} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF39} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hF3A} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF3D} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hF3E} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b011, 12'hF41} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b011, 12'hF42} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF43} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF45} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b011, 12'hF46} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF47} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF49} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b011, 12'hF4A} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF4B} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF4D} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b011, 12'hF4E} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF4F} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF51} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b011, 12'hF52} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF53} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF55} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b011, 12'hF56} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF57} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF59} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b011, 12'hF5A} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF5B} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF5D} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b011, 12'hF5E} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF5F} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF61} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b011, 12'hF62} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF63} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF65} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b011, 12'hF66} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF67} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF69} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b011, 12'hF6A} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF6B} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF6D} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b011, 12'hF6E} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF6F} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF71} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hF72} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF73} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF75} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hF76} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF77} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF79} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hF7A} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF7B} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF7D} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b011, 12'hF7E} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b011, 12'hF7F} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b011, 12'hF80} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b011, 12'hF84} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b011, 12'hF88} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b011, 12'hF8C} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b011, 12'hF90} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b011, 12'hF94} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b011, 12'hF98} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b011, 12'hF9C} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b011, 12'hFA0} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b011, 12'hFA4} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b011, 12'hFA8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b011, 12'hFAC} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b011, 12'hFB0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b011, 12'hFB4} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b011, 12'hFB8} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b011, 12'hFBC} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b011, 12'hFC0} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b011, 12'hFC4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b011, 12'hFC8} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b011, 12'hFCC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b011, 12'hFD0} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b011, 12'hFD4} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b011, 12'hFD8} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b011, 12'hFDC} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b011, 12'hFE0} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b011, 12'hFE4} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b011, 12'hFE8} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b011, 12'hFEC} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b011, 12'hFF0} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b011, 12'hFF4} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b011, 12'hFF8} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b011, 12'hFFC} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b100, 12'h001} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h004} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h005} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h008} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h009} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h00C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h00D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h010} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h011} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h014} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b100, 12'h015} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h018} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b100, 12'h019} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h01C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h01D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h020} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h021} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h024} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'h025} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h028} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h029} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h02C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h02D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h030} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h031} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h034} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h035} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h038} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h039} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h03C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h03D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h040} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h041} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h044} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b100, 12'h045} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h048} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b100, 12'h049} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h04C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b100, 12'h04D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h050} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b100, 12'h051} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h054} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b100, 12'h055} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h058} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b100, 12'h059} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h05C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b100, 12'h05D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h060} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b100, 12'h061} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h064} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b100, 12'h065} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h068} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h069} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h06C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b100, 12'h06D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h070} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h071} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h074} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b100, 12'h075} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h078} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b100, 12'h079} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h07C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'h07D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h080} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h081} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h084} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b100, 12'h085} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h088} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'h089} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h08C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b100, 12'h08D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h090} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b100, 12'h091} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h094} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b100, 12'h095} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h098} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b100, 12'h099} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h09C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b100, 12'h09D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0A0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b100, 12'h0A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0A4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'h0A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0A8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'h0A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0AC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b100, 12'h0AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0B0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h0B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0B4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h0B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0B8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h0B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0BC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h0BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0C0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h0C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0C4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b100, 12'h0C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0C8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b100, 12'h0C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0CC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b100, 12'h0CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0D0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b100, 12'h0D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0D4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b100, 12'h0D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0D8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b100, 12'h0D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0DC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b100, 12'h0DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0E0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b100, 12'h0E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0E4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b100, 12'h0E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0E8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b100, 12'h0E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0EC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b100, 12'h0ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0F0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b100, 12'h0F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0F4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b100, 12'h0F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b100, 12'h0F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h0FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b100, 12'h0FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h100} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h101} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h104} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b100, 12'h105} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h108} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b100, 12'h109} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h10C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b100, 12'h10D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h110} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b100, 12'h111} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h114} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b100, 12'h115} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h118} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b100, 12'h119} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h11C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b100, 12'h11D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h120} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b100, 12'h121} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h124} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b100, 12'h125} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h128} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b100, 12'h129} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h12C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b100, 12'h12D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h130} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b100, 12'h131} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h134} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b100, 12'h135} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h138} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b100, 12'h139} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h13C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'h13D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h140} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h141} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h144} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b100, 12'h145} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h148} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b100, 12'h149} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h14C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b100, 12'h14D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h150} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b100, 12'h151} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h154} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b100, 12'h155} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h158} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b100, 12'h159} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h15C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b100, 12'h15D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h160} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b100, 12'h161} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h164} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b100, 12'h165} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h168} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b100, 12'h169} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h16C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b100, 12'h16D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h170} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b100, 12'h171} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h174} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b100, 12'h175} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h178} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b100, 12'h179} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h17C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b100, 12'h17D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h180} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h181} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h184} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b100, 12'h185} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h188} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b100, 12'h189} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h18C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b100, 12'h18D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h190} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b100, 12'h191} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h194} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b100, 12'h195} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h198} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b100, 12'h199} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h19C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b100, 12'h19D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b100, 12'h1A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b100, 12'h1A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b100, 12'h1A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b100, 12'h1AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b100, 12'h1B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b100, 12'h1B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b100, 12'h1B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b100, 12'h1BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1C0} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b100, 12'h1C1} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b100, 12'h1C2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h1C4} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h1C5} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h1C6} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'h1C8} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b100, 12'h1C9} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b100, 12'h1CA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h1CB} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h1CC} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'h1CE} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b100, 12'h1CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h1D0} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b100, 12'h1D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1D4} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b100, 12'h1D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1D8} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b100, 12'h1D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1DC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b100, 12'h1E0} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b100, 12'h1E4} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h1E8} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h1EC} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h1F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b100, 12'h1F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h1F2} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b100, 12'h1F4} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b100, 12'h1F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h1F6} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b100, 12'h1F8} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b100, 12'h1FC} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b100, 12'h201} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h202} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h204} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b100, 12'h206} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h207} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h208} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'h209} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'h20E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h211} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h213} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h215} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h219} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h21B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h21D} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h21E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h220} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b100, 12'h222} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h224} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b100, 12'h226} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h227} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h228} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b100, 12'h229} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'h22E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h231} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h233} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h235} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h239} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h23B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h23E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h240} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h242} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h244} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b100, 12'h245} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b100, 12'h246} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b100, 12'h248} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b100, 12'h249} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b100, 12'h24A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h24D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h24E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h251} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b100, 12'h252} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b100, 12'h255} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h256} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h259} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'h25A} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b100, 12'h25D} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'h25E} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'h261} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h262} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h263} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h265} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b100, 12'h266} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'h269} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h26A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h26B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h26C} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h26D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h26F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h270} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b100, 12'h271} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b100, 12'h272} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h273} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h275} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h277} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h278} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h279} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h27B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h27C} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'h27D} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b100, 12'h281} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h283} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h285} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h289} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h28A} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h28B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h28D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h28E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h28F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h290} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h291} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h293} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h294} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b100, 12'h295} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b100, 12'h296} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h297} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h299} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h29B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h29C} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h2A0} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b100, 12'h2A1} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b100, 12'h2A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2A5} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h2A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2A9} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h2AD} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h2AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2B0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h2B1} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h2B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2B4} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b100, 12'h2B5} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'h2B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2B8} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'h2B9} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b100, 12'h2BA} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h2BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2BC} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'h2BD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'h2BE} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h2BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2C0} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'h2C1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h2C2} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'h2C4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b100, 12'h2C5} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h2C8} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'h2C9} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h2CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2CD} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2CE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h2CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2D4} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'h2D5} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h2D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2D9} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2DA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h2DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2DE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h2DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2E0} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'h2E1} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h2E2} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h2E4} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h2E5} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h2E6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2E8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h2E9} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h2EA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h2EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h2EC} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b100, 12'h2ED} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'h2F0} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b100, 12'h2F1} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h2F5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h2F6} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h2FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h2FE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h300} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h301} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h302} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h303} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h305} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h306} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b100, 12'h307} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h309} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h30D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h311} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h312} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'h313} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h314} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h315} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h319} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h31A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h31B} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'h321} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h322} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h323} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h324} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'h325} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h326} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h328} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h329} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h32A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h32B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h32C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b100, 12'h32D} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'h331} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h332} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h333} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h335} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h336} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h337} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h338} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b100, 12'h339} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b100, 12'h33B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h33C} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b100, 12'h33D} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h341} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h342} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h349} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h34A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h34C} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h34D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h34E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h34F} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h351} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h352} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b100, 12'h353} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h355} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h356} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h357} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h358} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h359} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h35D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h35E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h35F} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'h365} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h366} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h367} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h36A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h36B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h36D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h36E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h36F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h370} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h371} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h373} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h374} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h375} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h376} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h377} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h378} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h379} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h37A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h37C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b100, 12'h37D} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h37E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h37F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h381} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h382} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h383} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h386} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h389} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h38A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h38B} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h38C} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b100, 12'h38D} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b100, 12'h38E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h38F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h390} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h391} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h393} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h394} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b100, 12'h395} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h39B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h39C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h39D} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h39F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3A0} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b100, 12'h3A1} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b100, 12'h3A2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h3A5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h3A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3A9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h3AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3AC} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h3AE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h3B0} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b100, 12'h3B1} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b100, 12'h3B2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h3B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3B4} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'h3B5} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h3B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3B8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b100, 12'h3B9} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h3BA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h3BB} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h3BC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'h3BD} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h3BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3C0} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h3C1} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'h3C5} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h3C6} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h3C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3C9} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h3CA} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h3CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h3CE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h3CF} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h3D0} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b100, 12'h3D1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h3D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3D5} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h3D6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h3D7} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h3DD} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h3DE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h3DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3E0} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b100, 12'h3E1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h3E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3E4} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h3E5} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h3E6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h3E7} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h3E9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'h3ED} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h3EE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h3EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3F1} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h3F2} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h3F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h3F6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h3F7} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h3F8} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b100, 12'h3F9} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h3FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h3FD} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h3FE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h3FF} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h405} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h406} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h407} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h408} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b100, 12'h409} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h40B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h40D} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h40E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h40F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h411} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h413} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h414} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h416} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h418} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b100, 12'h419} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h41A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h41B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h41D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h41E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h420} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h421} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h422} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h423} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h425} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h426} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h427} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h428} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h429} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h42A} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'h42B} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h42C} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h430} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b100, 12'h431} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h433} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'h435} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b100, 12'h436} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h437} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h439} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'h43A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h43B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h43C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h43D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h43F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h440} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b100, 12'h441} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b100, 12'h442} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h443} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h445} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b100, 12'h447} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h449} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b100, 12'h44B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h44C} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b100, 12'h44D} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b100, 12'h450} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h453} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h454} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b100, 12'h455} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h458} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h459} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b100, 12'h45A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h45B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h45D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h45E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h461} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h463} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h464} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h465} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h466} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h467} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h468} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b100, 12'h469} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b100, 12'h46B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h46D} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h471} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h472} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h475} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h477} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h478} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h479} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h47A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h47B} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h47C} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b100, 12'h47D} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b100, 12'h47F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h480} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h481} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b100, 12'h484} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h486} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h487} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h488} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b100, 12'h489} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b100, 12'h48A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h48C} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h48D} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b100, 12'h48E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h48F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h490} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h491} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h493} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h494} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b100, 12'h495} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b100, 12'h496} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h497} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h499} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h49A} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h49C} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h49D} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h49E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h49F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h4A2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h4A3} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h4A5} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h4A6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h4A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4A9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h4AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h4AE} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h4B0} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4B1} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b100, 12'h4B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4B4} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h4B8} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b100, 12'h4B9} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h4BA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h4BB} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h4BD} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h4BE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h4BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4C1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h4C5} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h4C6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h4C7} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h4C8} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4C9} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h4CA} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h4CC} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h4D0} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b100, 12'h4D1} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h4D4} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h4D7} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'h4D8} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h4D9} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b100, 12'h4DA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h4DB} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h4DD} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h4DE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h4E0} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h4E1} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h4E2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h4E6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h4E7} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h4E9} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h4EA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h4EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4ED} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h4F4} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h4F5} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h4F6} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h4F8} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h4FC} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b100, 12'h4FD} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h4FE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h4FF} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h501} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h502} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h503} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h505} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h509} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h50A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h50B} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h50C} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h50D} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h50E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h510} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h514} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b100, 12'h515} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h518} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h51B} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'h51C} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h51D} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b100, 12'h51E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h51F} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h520} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h521} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h523} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h524} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b100, 12'h525} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h526} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h527} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h528} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h52A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h52C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h52E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h531} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h532} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h533} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h536} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h537} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h53A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h53D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h53E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h53F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h541} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'h542} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b100, 12'h544} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'h545} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h546} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h548} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h54A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h54B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h54C} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b100, 12'h54D} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b100, 12'h54E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h54F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h550} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b100, 12'h551} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'h554} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b100, 12'h555} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h557} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h559} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h55A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h55D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h55E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h55F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h561} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'h564} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b100, 12'h565} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h569} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h56D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h570} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b100, 12'h571} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'h574} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b100, 12'h575} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h57C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h57D} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'h57E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h57F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h580} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b100, 12'h581} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h582} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h583} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h585} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h586} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h589} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h58B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h58D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h58E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h58F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h590} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b100, 12'h591} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h592} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h594} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h595} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h596} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h59A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h59D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h59E} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'h5A0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h5A2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h5A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5A4} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b100, 12'h5A5} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h5A8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b100, 12'h5A9} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h5AA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5AC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h5AD} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h5AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5B0} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b100, 12'h5B1} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b100, 12'h5B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5B5} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h5B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5B8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h5B9} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h5BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5BC} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b100, 12'h5BD} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b100, 12'h5BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5C1} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h5C2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h5C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5C8} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b100, 12'h5C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h5CA} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b100, 12'h5CC} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h5CD} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h5CE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h5CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5D0} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b100, 12'h5D1} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'h5D5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h5D6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h5D7} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h5D8} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h5D9} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b100, 12'h5DA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h5DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5DC} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b100, 12'h5DD} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h5E0} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h5E1} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'h5E2} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b100, 12'h5E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h5E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h5EA} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h5EC} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h5ED} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h5EE} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h5EF} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h5F0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b100, 12'h5F1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h5F2} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b100, 12'h5F3} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h5F9} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h5FA} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b100, 12'h5FB} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h5FC} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h5FD} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h601} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h602} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'h603} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h605} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h606} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h609} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h60A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h60B} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h60D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h615} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h616} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h617} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h619} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'h61A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h61B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h61D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h61F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h620} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h622} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h624} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b100, 12'h625} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b100, 12'h626} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h627} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h628} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h629} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h62A} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b100, 12'h62B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h62D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h62F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h630} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h631} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h632} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h633} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h635} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h636} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b100, 12'h637} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h639} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h63A} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h63B} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h63C} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h63D} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h640} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h641} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h642} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h643} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h644} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b100, 12'h645} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h646} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h647} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h648} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h649} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h64B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h64C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b100, 12'h64D} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'h64E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h64F} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'h650} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h652} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h654} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h656} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h659} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h65A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h65B} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h65D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h65E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h65F} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'h660} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h661} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h662} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h664} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h666} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h668} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'h669} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b100, 12'h66A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h66B} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h66E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h66F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h670} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b100, 12'h671} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h672} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h676} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h679} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h67A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h67B} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h67D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h67E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h67F} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'h681} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h682} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h683} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h686} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h688} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'h689} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b100, 12'h68A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h68B} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h68C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h68D} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h68F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h690} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b100, 12'h691} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'h692} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h695} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h697} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h698} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b100, 12'h699} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h69A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h69C} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'h69D} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h69E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h69F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6A0} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b100, 12'h6A1} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h6A2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h6A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6A5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h6A6} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h6A9} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h6AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h6AE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h6B1} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h6B2} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h6B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6B5} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h6B6} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'h6B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6BE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h6BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6C0} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h6C1} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h6C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6C5} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h6C6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h6C7} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h6C9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h6CA} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h6CB} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h6CC} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h6D0} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b100, 12'h6D1} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b100, 12'h6D2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h6D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6D4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h6D5} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h6D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6D8} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b100, 12'h6D9} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b100, 12'h6DA} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'h6DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6DC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b100, 12'h6DE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6E0} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b100, 12'h6E1} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h6E2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h6E3} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h6E4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h6E5} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h6E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6E8} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b100, 12'h6E9} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h6EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6F0} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b100, 12'h6F1} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h6F2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h6F3} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h6F4} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b100, 12'h6F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h6F8} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b100, 12'h6F9} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h6FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h6FC} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h6FD} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h6FE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h6FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h700} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b100, 12'h701} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b100, 12'h702} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h703} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h705} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h707} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h708} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h70B} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'h70C} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b100, 12'h70D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h714} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'h715} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h717} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h718} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'h719} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h71C} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b100, 12'h71D} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b100, 12'h721} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h724} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h725} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h726} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h727} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h728} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h72A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h72C} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b100, 12'h72D} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b100, 12'h72E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h730} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b100, 12'h731} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h732} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h733} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h735} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h736} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h737} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h739} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h73A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h73B} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h73C} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h73D} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h73E} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'h73F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h740} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h741} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h743} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h745} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h749} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h74A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h74B} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h74D} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h74E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h74F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h750} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'h751} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h752} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h755} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b100, 12'h757} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h758} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h75C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b100, 12'h75D} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'h760} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'h761} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h763} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h764} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b100, 12'h765} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h766} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h767} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h768} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h769} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h76A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h76B} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h76C} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b100, 12'h76D} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'h76F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h770} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b100, 12'h771} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h774} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h775} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h776} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'h778} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'h779} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b100, 12'h77A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h77C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h77D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'h77F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h780} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'h781} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h782} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h783} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h784} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'h785} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h788} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'h789} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b100, 12'h78A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h78C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h78F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h790} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h791} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h794} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h795} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h796} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b100, 12'h798} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b100, 12'h799} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h79A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h79B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h79D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h79E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h79F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7A1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h7A2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7A4} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b100, 12'h7A5} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b100, 12'h7A6} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'h7A7} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h7A9} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h7AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7AC} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b100, 12'h7AD} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h7AE} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'h7AF} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h7B0} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h7B4} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b100, 12'h7B5} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h7B6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h7B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7B8} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b100, 12'h7B9} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h7BA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h7BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7BC} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b100, 12'h7BD} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h7BE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h7BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7C0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b100, 12'h7C1} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b100, 12'h7C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7C4} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h7C5} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h7C8} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b100, 12'h7CA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7CC} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b100, 12'h7CD} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b100, 12'h7CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7D0} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b100, 12'h7D2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7D4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b100, 12'h7D5} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b100, 12'h7D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7D8} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h7DA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7DC} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b100, 12'h7DD} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b100, 12'h7DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7E0} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h7E2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7E4} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b100, 12'h7E5} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b100, 12'h7E7} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h7E8} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'h7EA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7EC} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7ED} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h7EE} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'h7EF} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h7F4} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h7F5} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h7F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h7F9} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h7FA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h7FB} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h7FC} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h7FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h7FE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h7FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h800} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h803} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h804} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h805} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b100, 12'h806} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h807} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h808} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'h80C} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'h80D} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h80E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h814} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h815} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h816} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h817} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h81C} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h81F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h820} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h821} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h822} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h823} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h824} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h825} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h827} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h828} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'h829} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h82A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h82B} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h82C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h82F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h830} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h831} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h832} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h834} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h835} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h836} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h837} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h838} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b100, 12'h839} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h83A} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'h83C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h83D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h83E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h83F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h840} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b100, 12'h841} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'h842} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h843} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'h844} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b100, 12'h845} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h848} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b100, 12'h849} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b100, 12'h84B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h84C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h84E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h84F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h850} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b100, 12'h851} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b100, 12'h853} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h854} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b100, 12'h855} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h856} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h857} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h858} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h859} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'h85B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h85C} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b100, 12'h85D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h864} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h865} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h867} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h868} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h869} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'h86A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h86B} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'h86C} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h86D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h876} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h878} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b100, 12'h87A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h881} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h882} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h883} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h885} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h886} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h887} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h888} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'h889} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b100, 12'h88B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h88C} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b100, 12'h88D} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'h88E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h895} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h896} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b100, 12'h897} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h898} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h899} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b100, 12'h89B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h89D} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b100, 12'h89E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h89F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h8A0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h8A1} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h8A2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h8A4} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h8A5} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h8A6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8A7} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h8A8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h8A9} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h8AA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8AC} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h8AD} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b100, 12'h8AE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8B1} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h8B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h8B5} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h8B6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8B9} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'h8BA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8BD} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b100, 12'h8BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h8C2} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b100, 12'h8C4} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b100, 12'h8C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h8C8} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b100, 12'h8C9} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b100, 12'h8CA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8CB} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h8CC} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b100, 12'h8CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h8CE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h8CF} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h8D1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h8D2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h8D3} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h8D5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h8D6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8D7} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h8D8} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h8D9} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h8DA} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'h8DB} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h8DC} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h8DD} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h8DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h8E1} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h8E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h8E6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h8E7} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h8E9} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'h8EA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h8EC} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'h8ED} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h8EE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h8F0} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b100, 12'h8F1} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b100, 12'h8F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h8F4} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h8F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h8F8} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h8F9} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b100, 12'h8FC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'h900} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h901} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h904} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'h905} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h906} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h907} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h908} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h909} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b100, 12'h90B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h90C} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h90D} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h910} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h914} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h915} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b100, 12'h917} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h918} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'h91B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h91C} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h91D} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b100, 12'h920} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'h921} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h922} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h928} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h929} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'h92A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'h92B} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'h930} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h933} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h934} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h935} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h936} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h937} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h938} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h939} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h93B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h93D} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h93E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h93F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'h940} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'h941} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b100, 12'h942} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h944} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'h945} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h946} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h948} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h94A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h94B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h94C} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b100, 12'h94D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h94E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h94F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h950} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b100, 12'h951} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h954} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b100, 12'h955} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h957} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h959} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'h95C} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b100, 12'h95D} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h961} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h964} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h965} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'h966} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h967} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h968} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b100, 12'h96A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h96B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h970} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b100, 12'h971} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h972} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b100, 12'h974} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b100, 12'h975} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h976} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h979} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'h97A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h97B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h97D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h981} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'h985} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h98C} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'h98D} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b100, 12'h98E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'h991} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b100, 12'h992} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h995} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'h996} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b100, 12'h998} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'h999} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h99A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h99B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h99E} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'h99F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9A6} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b100, 12'h9AD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'h9AE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'h9B0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'h9B1} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h9B2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h9B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9B4} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b100, 12'h9B5} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'h9B7} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'h9B8} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b100, 12'h9B9} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'h9BC} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'h9BD} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b100, 12'h9BE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h9C0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h9C1} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'h9C2} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'h9C6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h9C7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9C9} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'h9CA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h9CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9CD} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b100, 12'h9CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9D5} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h9D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9D8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h9D9} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'h9DA} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h9DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9DC} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b100, 12'h9DD} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b100, 12'h9DE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'h9DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9E1} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h9E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9E4} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'h9E5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h9E6} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'h9E7} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'h9E8} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'h9E9} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'h9EC} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b100, 12'h9ED} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'h9EE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'h9F0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'h9F1} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'h9F2} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'h9F4} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b100, 12'h9F5} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'h9F6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9F8} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b100, 12'h9F9} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b100, 12'h9FA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'h9FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA05} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hA06} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'hA08} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'hA09} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hA0A} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hA0B} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hA0D} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'hA0E} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b100, 12'hA0F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hA11} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hA12} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hA13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA14} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hA15} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'hA19} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hA1A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hA1B} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'hA1D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hA1E} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'hA20} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b100, 12'hA21} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b100, 12'hA22} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hA23} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hA24} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b100, 12'hA25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hA26} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA29} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hA2D} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'hA2E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hA2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA30} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b100, 12'hA31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hA34} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'hA35} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b100, 12'hA36} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hA38} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'hA39} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hA3A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hA3C} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'hA3E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hA3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA41} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA44} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'hA45} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hA46} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hA47} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hA48} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b100, 12'hA49} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hA4B} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hA4D} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hA50} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b100, 12'hA51} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b100, 12'hA53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA54} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hA55} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hA57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA58} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'hA59} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hA5A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hA5B} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hA5C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hA5D} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hA5E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA60} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b100, 12'hA61} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'hA65} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hA66} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hA67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA6A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA6D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hA6E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hA6F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hA71} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b100, 12'hA72} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hA74} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hA75} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hA77} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA78} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b100, 12'hA79} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b100, 12'hA7A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA7D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'hA80} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hA81} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'hA82} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hA83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA84} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hA85} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'hA86} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hA87} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA88} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hA89} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'hA8A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hA8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA8D} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'hA8E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hA8F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hA90} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hA91} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hA92} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hA93} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hA94} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b100, 12'hA95} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b100, 12'hA98} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hA99} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'hA9A} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b100, 12'hA9D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hA9F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAA1} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hAA3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAA4} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hAA5} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b100, 12'hAA6} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hAA7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAA9} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hAAA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hAAB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAAD} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hAAE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAAF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAB0} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hAB1} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b100, 12'hAB2} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hAB3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAB5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hAB6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hAB7} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hAB9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hABD} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b100, 12'hABF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAC1} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'hAC2} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hAC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAC5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hAC6} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hAC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAC9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hACA} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b100, 12'hACB} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hACD} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b100, 12'hACE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hACF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAD0} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b100, 12'hAD3} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'hAD5} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b100, 12'hAD9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hADA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hADB} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hADD} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b100, 12'hADE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hADF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAE0} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'hAE1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hAE3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAE4} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hAE5} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b100, 12'hAE6} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hAE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAE8} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'hAE9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hAEA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hAEB} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hAEC} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'hAED} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b100, 12'hAEE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hAEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAF0} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b100, 12'hAF1} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hAF3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAF4} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hAF5} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b100, 12'hAF9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hAFA} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hAFB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hAFC} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b100, 12'hAFD} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hAFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB00} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'hB01} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'hB05} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hB07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB08} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hB09} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'hB0A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hB0B} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hB10} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b100, 12'hB11} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'hB12} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hB13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB15} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hB16} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hB17} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hB18} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hB1B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB1C} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b100, 12'hB1D} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'hB21} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b100, 12'hB22} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hB23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB25} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hB26} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hB28} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hB2A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hB2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB2C} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b100, 12'hB2D} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b100, 12'hB2E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hB2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB30} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b100, 12'hB31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hB32} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB33} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB34} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hB35} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hB37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB38} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b100, 12'hB39} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b100, 12'hB3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB3C} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b100, 12'hB3D} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'hB3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB40} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b100, 12'hB41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hB44} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'hB46} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB47} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB48} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hB49} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hB4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB4C} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b100, 12'hB4D} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hB4E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hB4F} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hB51} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hB54} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b100, 12'hB55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hB5A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB62} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hB65} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'hB66} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hB68} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hB69} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hB6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB6C} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b100, 12'hB6D} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hB6E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hB6F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hB70} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'hB71} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'hB73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB74} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b100, 12'hB75} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b100, 12'hB76} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hB77} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB79} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'hB7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB7E} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b100, 12'hB80} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hB81} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hB83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB84} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b100, 12'hB85} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hB86} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hB87} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hB88} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b100, 12'hB89} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hB8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB8D} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b100, 12'hB8E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hB8F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB90} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b100, 12'hB91} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b100, 12'hB93} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB97} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hB98} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hB99} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'hB9A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hB9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hB9C} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b100, 12'hB9D} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b100, 12'hB9E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hBA0} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'hBA1} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b100, 12'hBA2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hBA5} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hBA7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hBA9} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'hBAA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hBAD} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hBAE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hBB1} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hBB3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hBB6} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b100, 12'hBB8} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b100, 12'hBB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hBBC} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b100, 12'hBBD} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'hBBE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hBBF} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'hBC0} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'hBC4} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b100, 12'hBC5} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hBC6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hBC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hBC9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hBCB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hBD1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hBD2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'hBD4} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'hBD5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hBD6} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hBD7} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hBD9} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'hBDA} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b100, 12'hBDB} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hBDC} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hBDD} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'hBE0} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b100, 12'hBE1} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'hBE2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hBE3} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hBE5} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'hBE6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hBE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hBE9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hBEA} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hBEB} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hBED} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hBEE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hBF1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hBF2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hBF3} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hBF5} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hBF6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hBF7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hBF8} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b100, 12'hBF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hBFA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hBFB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hBFC} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b100, 12'hBFD} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b100, 12'hBFE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hC00} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'hC01} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b100, 12'hC02} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hC03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC06} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hC07} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC09} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hC0A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC0B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC0C} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hC0D} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b100, 12'hC0E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hC0F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC10} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hC11} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b100, 12'hC13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC15} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'hC19} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'hC1B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC1D} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hC1F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC20} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hC21} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b100, 12'hC22} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hC23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC24} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hC25} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'hC26} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hC27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC29} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'hC2A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hC2B} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hC2F} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'hC31} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hC34} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hC35} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hC36} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hC37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC38} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b100, 12'hC39} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'hC3D} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hC3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC41} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b100, 12'hC42} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hC45} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hC47} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC49} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hC4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC4D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hC4E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hC4F} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hC51} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hC52} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hC54} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hC55} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hC56} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hC57} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hC59} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b100, 12'hC5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC5D} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b100, 12'hC5E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hC5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC65} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hC66} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hC67} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hC68} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hC69} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'hC6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC6C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b100, 12'hC6D} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b100, 12'hC6E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hC6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC70} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b100, 12'hC73} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'hC75} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b100, 12'hC81} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hC82} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hC83} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hC84} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'hC85} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'hC87} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC88} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hC89} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b100, 12'hC8A} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hC8C} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hC8D} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'hC8F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC90} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b100, 12'hC91} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hC95} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'hC96} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hC97} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hC99} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hC9C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hCA0} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'hCA1} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hCA2} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hCA4} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b100, 12'hCA7} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'hCA8} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hCA9} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hCAC} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'hCAD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hCAE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hCAF} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hCB0} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b100, 12'hCB1} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hCB3} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b100, 12'hCB4} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hCB5} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b100, 12'hCB9} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'hCBA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hCBC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hCBE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hCBF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hCC0} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'hCC1} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b100, 12'hCC4} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b100, 12'hCC5} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'hCC6} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hCC8} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b100, 12'hCC9} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hCCB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hCCC} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b100, 12'hCCD} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hCCE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hCD1} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'hCD3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hCD5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hCD6} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b100, 12'hCD7} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hCD8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hCD9} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hCDB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hCDD} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b100, 12'hCDF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hCE4} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b100, 12'hCE5} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'hCE6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hCE7} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hCE8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hCE9} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hCEB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hCEC} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b100, 12'hCED} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hCEE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hCEF} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hCF0} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hCF1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hCF2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hCF4} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hCF6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hCF8} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hCF9} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b100, 12'hCFB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hCFC} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'hCFD} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hCFE} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hCFF} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hD00} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hD01} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hD02} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD04} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hD05} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b100, 12'hD0D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hD0E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hD0F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hD10} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hD11} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hD12} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hD13} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD14} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'hD15} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'hD18} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hD19} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'hD1A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hD1B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD1C} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b100, 12'hD1D} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hD1E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hD20} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'hD21} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hD23} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD24} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b100, 12'hD25} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hD28} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b100, 12'hD29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hD2D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hD2E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hD2F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hD30} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hD31} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'hD32} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hD33} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hD34} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hD35} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'hD37} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD39} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hD3D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hD3E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hD3F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hD40} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hD43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD44} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'hD45} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b100, 12'hD46} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hD48} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'hD49} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b100, 12'hD4A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hD4D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hD4E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD52} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD55} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hD56} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hD58} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hD5A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hD5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD5C} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'hD5D} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hD5E} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hD5F} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hD60} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hD61} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hD62} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD63} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD64} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hD65} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b100, 12'hD68} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b100, 12'hD69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hD6C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'hD6D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'hD6E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hD70} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hD71} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hD72} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hD73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD74} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b100, 12'hD75} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hD76} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hD77} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD78} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'hD79} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b100, 12'hD7A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hD7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD7C} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b100, 12'hD7D} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hD7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD81} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hD82} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hD83} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD84} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b100, 12'hD85} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b100, 12'hD86} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hD89} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hD8A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hD8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hD8D} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'hD8E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hD91} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hD94} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b100, 12'hD95} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'hD99} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'hD9C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hD9D} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hD9E} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'hD9F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDA0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b100, 12'hDA2} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'hDA3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDA8} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b100, 12'hDA9} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hDAA} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b100, 12'hDAC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b100, 12'hDAD} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'hDAE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDB1} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hDB2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDB3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDB5} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'hDB6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hDB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDBC} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hDBD} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b100, 12'hDBE} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'hDC1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hDC2} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hDC6} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'hDC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDCE} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b100, 12'hDD5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hDD6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hDD9} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'hDDA} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b100, 12'hDDC} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b100, 12'hDDD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hDDE} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hDE0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hDE1} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'hDE2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hDE3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDE4} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b100, 12'hDE5} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b100, 12'hDE8} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'hDE9} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hDEA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDEB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDEC} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b100, 12'hDED} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'hDF0} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'hDF1} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hDF2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDF3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDF5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hDF6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hDF7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hDF8} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b100, 12'hDF9} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'hDFC} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b100, 12'hDFD} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b100, 12'hE01} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hE02} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hE09} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hE0A} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b100, 12'hE0C} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'hE0D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hE0E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hE0F} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hE11} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b100, 12'hE12} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b100, 12'hE13} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hE15} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hE16} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hE17} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hE18} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'hE19} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hE1A} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'hE1C} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b100, 12'hE1D} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b100, 12'hE20} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b100, 12'hE22} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE26} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE28} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b100, 12'hE29} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'hE2A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hE2B} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hE2C} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'hE2D} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hE2E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE2F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE30} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hE31} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b100, 12'hE33} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE34} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hE35} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'hE36} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'hE37} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'hE3A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hE3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE3D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'hE3E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE3F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE40} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b100, 12'hE42} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE45} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hE46} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hE47} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE49} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hE4A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hE4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE4C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hE4D} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b100, 12'hE4E} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hE4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE52} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hE53} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE54} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b100, 12'hE55} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hE56} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hE58} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hE5A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hE5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE5C} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b100, 12'hE5D} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'hE5E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE5F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE60} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b100, 12'hE64} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b100, 12'hE65} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b100, 12'hE67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE68} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b100, 12'hE69} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hE6A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hE6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE6C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hE6E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hE70} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b100, 12'hE71} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hE74} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b100, 12'hE76} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE78} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b100, 12'hE79} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hE7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE7C} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b100, 12'hE7D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hE7E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hE7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE80} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hE82} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hE84} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b100, 12'hE85} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'hE86} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hE88} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b100, 12'hE8A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE8C} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b100, 12'hE8D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hE8E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE90} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b100, 12'hE91} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'hE92} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hE93} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE95} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hE96} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hE98} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b100, 12'hE99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hE9A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hE9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hE9C} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hE9E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEA0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b100, 12'hEA1} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b100, 12'hEA2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEA3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEA4} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hEA6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEA8} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b100, 12'hEA9} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hEAC} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b100, 12'hEAD} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hEB2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hEB4} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b100, 12'hEB5} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b100, 12'hEB6} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hEB9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hEBA} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hEBC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hEBE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hEBF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEC0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b100, 12'hEC1} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b100, 12'hEC2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hEC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEC4} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hEC8} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b100, 12'hEC9} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hECE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hECF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hED1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hED2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hED3} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hED5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hED6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hED7} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hED9} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hEDA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b100, 12'hEDB} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b100, 12'hEDC} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b100, 12'hEDD} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b100, 12'hEE0} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hEE1} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hEE2} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hEE5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hEE6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEE9} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'hEEB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEEC} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b100, 12'hEED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hEEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEF0} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'hEF2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEF3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEF4} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b100, 12'hEF5} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b100, 12'hEF6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hEF7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hEF8} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'hEFC} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b100, 12'hEFD} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hEFE} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'hEFF} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b100, 12'hF00} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b100, 12'hF01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hF02} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF03} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF05} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hF06} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hF08} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b100, 12'hF0A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF0E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF11} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hF12} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hF13} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b100, 12'hF14} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b100, 12'hF16} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF17} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF18} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b100, 12'hF1C} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b100, 12'hF1D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hF1E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hF21} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b100, 12'hF22} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b100, 12'hF23} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hF25} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b100, 12'hF26} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hF27} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF28} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hF29} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b100, 12'hF2A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hF2B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF2C} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b100, 12'hF2E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF30} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b100, 12'hF31} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b100, 12'hF32} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hF34} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b100, 12'hF36} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF38} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b100, 12'hF39} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hF3A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hF3B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF3C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hF3E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF40} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b100, 12'hF41} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hF42} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hF43} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF45} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hF46} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hF48} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hF4A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hF4B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF4C} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b100, 12'hF4D} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b100, 12'hF4F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF50} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hF52} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF54} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b100, 12'hF55} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hF57} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF58} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b100, 12'hF59} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'hF5B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF5D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hF5E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hF60} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'hF61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hF62} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF63} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF64} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hF65} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hF67} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF68} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b100, 12'hF69} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hF6B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF6D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hF6E} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hF6F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF70} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b100, 12'hF71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hF72} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF73} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF75} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b100, 12'hF76} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hF78} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hF79} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hF7A} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b100, 12'hF7B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF7C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hF7D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'hF7F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF80} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hF81} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b100, 12'hF84} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b100, 12'hF85} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b100, 12'hF86} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b100, 12'hF87} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hF88} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b100, 12'hF89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hF8A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hF8B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF8D} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b100, 12'hF8E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b100, 12'hF8F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF91} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hF92} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF93} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF94} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hF95} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'hF97} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF98} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hF99} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b100, 12'hF9A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF9B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF9C} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b100, 12'hF9D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'hF9E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hF9F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFA0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b100, 12'hFA1} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b100, 12'hFA2} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b100, 12'hFA4} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b100, 12'hFA6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFA8} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hFAA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFAC} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b100, 12'hFAD} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b100, 12'hFAE} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hFB0} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b100, 12'hFB1} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b100, 12'hFB2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hFB4} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hFB5} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b100, 12'hFB6} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hFB7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFB8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b100, 12'hFB9} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b100, 12'hFBA} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b100, 12'hFBB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFBC} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hFBD} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b100, 12'hFBE} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b100, 12'hFBF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFC1} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hFC2} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b100, 12'hFC3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFC4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b100, 12'hFC5} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b100, 12'hFC6} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hFC7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFC8} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b100, 12'hFC9} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b100, 12'hFCB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFCC} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b100, 12'hFCD} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b100, 12'hFCE} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b100, 12'hFCF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFD2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFD4} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b100, 12'hFD6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hFD8} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b100, 12'hFD9} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b100, 12'hFDC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b100, 12'hFDD} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b100, 12'hFDE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b100, 12'hFE0} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b100, 12'hFE1} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b100, 12'hFE5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b100, 12'hFE6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hFE7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFE9} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b100, 12'hFEA} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hFED} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hFEE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b100, 12'hFEF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFF0} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b100, 12'hFF1} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b100, 12'hFF3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFF5} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b100, 12'hFF6} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b100, 12'hFF7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b100, 12'hFF9} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b100, 12'hFFC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b100, 12'hFFD} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b100, 12'hFFF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h000} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h001} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h002} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h003} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h005} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h009} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h00A} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b101, 12'h00B} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h00C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h00D} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h00F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h010} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b101, 12'h011} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h012} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h013} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h014} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h018} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h019} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h01A} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b101, 12'h01B} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h01C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h01D} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h01E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h01F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h020} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b101, 12'h021} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h024} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b101, 12'h025} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h026} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h027} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h028} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b101, 12'h02A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h02B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h02D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h02E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h02F} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h030} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b101, 12'h034} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h035} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b101, 12'h037} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h038} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b101, 12'h039} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b101, 12'h03C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b101, 12'h03D} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b101, 12'h03E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h040} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h044} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b101, 12'h045} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b101, 12'h046} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h049} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b101, 12'h04B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h04D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h04E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h04F} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'h051} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'h055} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h057} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h058} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b101, 12'h059} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'h05A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h05B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h05D} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h060} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h061} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h062} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h063} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h064} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h065} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b101, 12'h066} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h067} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h068} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b101, 12'h069} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b101, 12'h06A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h06B} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b101, 12'h06C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h06D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b101, 12'h06E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h06F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h070} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h071} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h072} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h073} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'h074} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h075} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h076} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h078} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b101, 12'h079} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b101, 12'h07A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h07C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h07D} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h07E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h07F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h081} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h082} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h083} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h085} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h086} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h087} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h089} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h08A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h08D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h08E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h091} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h093} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h094} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h095} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h096} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b101, 12'h099} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b101, 12'h09A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h09D} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h09E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h09F} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h0A0} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b101, 12'h0A1} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h0A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0A5} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b101, 12'h0A6} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h0AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h0AE} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b101, 12'h0AF} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h0B0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h0B1} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h0B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0B5} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b101, 12'h0B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0BC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h0BD} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b101, 12'h0BE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h0BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0C0} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b101, 12'h0C1} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'h0C2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0C5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h0C6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h0C7} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b101, 12'h0C8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h0C9} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h0CC} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b101, 12'h0CD} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h0D0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h0D1} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b101, 12'h0D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0D5} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h0D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0D8} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h0D9} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b101, 12'h0DA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h0DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0DD} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b101, 12'h0DE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h0DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0E0} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b101, 12'h0E1} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b101, 12'h0E2} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h0E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0E5} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b101, 12'h0E6} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h0E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0E9} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'h0EA} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h0EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0EC} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h0ED} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b101, 12'h0EE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h0EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0F0} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b101, 12'h0F1} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'h0F2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0F5} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h0F8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h0F9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h0FA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h0FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h0FC} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b101, 12'h0FD} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b101, 12'h0FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h101} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h102} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h103} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b101, 12'h104} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b101, 12'h105} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b101, 12'h106} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h107} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h108} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h109} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h10B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h10C} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b101, 12'h10D} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h10E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h112} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h113} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h115} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h116} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h118} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b101, 12'h11A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h11B} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b101, 12'h11C} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b101, 12'h11D} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'h11E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h11F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h121} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b101, 12'h123} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h124} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h125} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b101, 12'h127} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h128} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h129} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h12A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h12B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h12C} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b101, 12'h12D} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'h12E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h12F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h132} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h133} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h134} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h138} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b101, 12'h139} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b101, 12'h13A} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h13B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h13C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h13D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h13F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h140} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b101, 12'h141} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b101, 12'h144} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b101, 12'h145} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h146} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h147} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h14A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h14B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h14C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h14D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h14E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h150} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h151} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b101, 12'h152} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h153} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h154} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h155} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b101, 12'h156} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h158} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h159} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h15A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h15B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h15C} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b101, 12'h15D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h15E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h15F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h160} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b101, 12'h161} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b101, 12'h162} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h163} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h164} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b101, 12'h165} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h167} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h169} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h16A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h16B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h16D} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b101, 12'h16E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h171} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h174} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b101, 12'h175} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b101, 12'h178} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b101, 12'h179} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b101, 12'h17D} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h17E} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h17F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h180} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b101, 12'h181} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b101, 12'h182} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h184} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h185} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b101, 12'h186} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b101, 12'h187} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h188} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b101, 12'h18A} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b101, 12'h18B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h190} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b101, 12'h191} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h192} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b101, 12'h194} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b101, 12'h195} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b101, 12'h196} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h199} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b101, 12'h19A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h19B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h19C} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h19D} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b101, 12'h19F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h1A1} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b101, 12'h1A2} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b101, 12'h1A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h1A4} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b101, 12'h1A5} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b101, 12'h1A6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h1A7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h1AA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h1AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h1AD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h1AE} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b101, 12'h1AF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h1B6} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b101, 12'h1B9} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h1BA} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h1BC} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h1BD} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b101, 12'h1BE} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h1BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h1C0} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b101, 12'h1C1} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'h1C5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h1C6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h1C7} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h1C8} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h1C9} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b101, 12'h1CA} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b101, 12'h1CC} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h1CD} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b101, 12'h1CE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h1CF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h1D0} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b101, 12'h1D1} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b101, 12'h1D2} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h1D4} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h1D5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h1D6} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h1D8} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b101, 12'h1D9} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b101, 12'h1DD} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h1DE} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h1E5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h1E6} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b101, 12'h1E8} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h1E9} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h1EA} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h1EB} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h1ED} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b101, 12'h1EE} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b101, 12'h1EF} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h1F0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h1F1} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b101, 12'h1F2} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b101, 12'h1F5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h1F6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h1F7} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'h1FD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h1FE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h1FF} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h200} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b101, 12'h201} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h202} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h203} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h204} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h205} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h207} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h208} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b101, 12'h209} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b101, 12'h20A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h20B} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b101, 12'h20C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h20E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h211} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h214} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b101, 12'h215} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b101, 12'h216} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h217} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h21A} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h21B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h21E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h221} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b101, 12'h223} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h224} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h225} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h226} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h227} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h228} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b101, 12'h229} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b101, 12'h22B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h22C} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b101, 12'h22D} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b101, 12'h22E} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h230} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b101, 12'h231} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h234} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h235} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b101, 12'h237} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h238} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b101, 12'h239} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b101, 12'h23B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h23C} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b101, 12'h23D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h23E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h23F} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'h240} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b101, 12'h241} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b101, 12'h243} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h244} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b101, 12'h245} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b101, 12'h248} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h249} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h24A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h24D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h24E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h24F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h250} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h251} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b101, 12'h252} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h253} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h255} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b101, 12'h256} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h258} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h25A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h25B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h25C} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b101, 12'h25D} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b101, 12'h25E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h25F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h261} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h262} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h263} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h264} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h265} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h267} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h268} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b101, 12'h269} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b101, 12'h26A} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h26B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h26D} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h26F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h270} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b101, 12'h271} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h276} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h277} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h279} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h27A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h27D} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h281} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b101, 12'h282} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h283} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h284} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h286} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h287} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h288} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b101, 12'h289} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b101, 12'h28A} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h28B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h28C} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b101, 12'h290} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b101, 12'h291} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h294} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h299} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b101, 12'h29A} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h29B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h29D} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h29F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2A0} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h2A2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2A4} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h2A5} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b101, 12'h2A8} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b101, 12'h2A9} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b101, 12'h2AA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h2AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2AC} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h2AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h2B0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h2B4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b101, 12'h2B5} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'h2B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2B9} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'h2BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2BC} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b101, 12'h2BD} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b101, 12'h2BE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2BF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2C0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h2C1} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h2C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2C4} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b101, 12'h2C5} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h2C8} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b101, 12'h2C9} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b101, 12'h2CA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2CC} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b101, 12'h2CD} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h2CE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2D0} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b101, 12'h2D1} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b101, 12'h2D2} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2D5} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h2D6} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2D8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h2DC} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b101, 12'h2DD} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b101, 12'h2DE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2DF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2E1} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h2E2} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h2E5} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h2E6} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b101, 12'h2E7} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h2E8} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h2E9} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b101, 12'h2EA} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b101, 12'h2EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2EC} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h2EE} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2F0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h2F1} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b101, 12'h2F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2F4} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b101, 12'h2F5} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b101, 12'h2F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h2F9} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h2FC} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b101, 12'h2FD} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b101, 12'h301} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h305} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h306} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h309} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h30A} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b101, 12'h30B} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h30D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b101, 12'h30F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h310} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h312} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h313} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h314} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b101, 12'h315} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b101, 12'h317} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h318} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b101, 12'h319} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h31C} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h31D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b101, 12'h31E} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h31F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h320} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b101, 12'h321} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b101, 12'h322} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b101, 12'h325} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b101, 12'h326} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h327} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h328} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h329} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h32B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h32C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b101, 12'h32D} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b101, 12'h32F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h330} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h331} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h332} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h333} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h335} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b101, 12'h337} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h339} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h33B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h340} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h341} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b101, 12'h342} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h344} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b101, 12'h345} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b101, 12'h346} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h347} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h34A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h34D} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h34E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h350} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h352} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h354} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b101, 12'h355} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b101, 12'h35A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h360} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h361} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h362} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h363} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h364} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h365} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b101, 12'h367} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h369} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h36A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h36B} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h36C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h36E} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h370} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h371} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b101, 12'h374} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b101, 12'h375} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b101, 12'h376} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h377} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h378} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b101, 12'h379} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h37A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h37C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h37D} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b101, 12'h37F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h380} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b101, 12'h381} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b101, 12'h382} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h385} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b101, 12'h387} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h389} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h38A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h38B} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'h38C} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b101, 12'h38D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h38F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h395} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'h398} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b101, 12'h399} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b101, 12'h39A} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h39B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h39D} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b101, 12'h39F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3A1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h3A2} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h3A5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h3A6} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h3A7} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h3A8} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h3A9} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h3AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3AC} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b101, 12'h3AD} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b101, 12'h3AE} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h3AF} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b101, 12'h3B0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h3B1} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'h3B3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3B4} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b101, 12'h3B5} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b101, 12'h3B7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3B8} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b101, 12'h3B9} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h3BA} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h3BB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3BC} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b101, 12'h3BD} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b101, 12'h3BE} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h3C1} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b101, 12'h3C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3C4} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b101, 12'h3C5} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h3C6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h3C7} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'h3C8} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b101, 12'h3C9} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b101, 12'h3CB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3CC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b101, 12'h3CD} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b101, 12'h3D1} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b101, 12'h3D2} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h3D4} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b101, 12'h3D5} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b101, 12'h3D8} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h3DA} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h3DB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3DC} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b101, 12'h3DD} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'h3E1} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h3E2} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h3E4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h3E6} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h3E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3E8} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b101, 12'h3E9} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h3EA} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h3EC} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h3EE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h3EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h3F0} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h3F1} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b101, 12'h3F5} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h3F6} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b101, 12'h3F8} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h3FC} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h3FD} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'h3FE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h3FF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h400} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h401} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h404} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b101, 12'h405} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h406} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h40A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h40B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h411} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h412} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h415} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h418} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b101, 12'h419} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b101, 12'h41A} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h41B} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h422} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h423} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h424} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h425} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h428} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b101, 12'h429} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h42A} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h42E} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h42F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h434} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h435} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h436} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h438} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b101, 12'h43C} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b101, 12'h43D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h43E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h43F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h441} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h442} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h444} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b101, 12'h446} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h447} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h448} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b101, 12'h449} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h44D} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h44E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h450} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h451} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h452} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h458} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b101, 12'h459} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h45B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h45C} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b101, 12'h45D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h460} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h461} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b101, 12'h462} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h465} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b101, 12'h466} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h468} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b101, 12'h469} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b101, 12'h46A} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h46B} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b101, 12'h46C} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h46D} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b101, 12'h46E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h46F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h470} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h471} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h472} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h473} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'h474} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h475} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h478} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h479} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h47A} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h47E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h47F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h480} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h482} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h484} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h485} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h488} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h48C} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b101, 12'h48D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h48E} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h48F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h494} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h495} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h496} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h499} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h49A} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h49B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h49C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h49D} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h49E} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h49F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4A1} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h4A2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h4A3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4A5} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h4A6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h4A9} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h4AB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4AE} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b101, 12'h4B0} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b101, 12'h4B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h4B4} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b101, 12'h4B5} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b101, 12'h4B6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h4B7} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b101, 12'h4B9} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b101, 12'h4BA} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h4BD} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h4BE} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h4BF} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h4C0} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b101, 12'h4C1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h4C3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4C5} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b101, 12'h4C6} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h4CD} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h4CE} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b101, 12'h4CF} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h4D0} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h4D1} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h4D3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4D5} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b101, 12'h4D7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4DD} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b101, 12'h4DE} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h4E1} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b101, 12'h4E2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h4E3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4E4} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h4E5} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b101, 12'h4E7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4E8} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b101, 12'h4E9} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b101, 12'h4EA} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h4EB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4EC} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b101, 12'h4ED} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b101, 12'h4EE} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h4EF} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4F1} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'h4F2} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h4F3} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4F4} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h4F5} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b101, 12'h4F6} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h4F7} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4F8} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b101, 12'h4F9} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b101, 12'h4FA} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h4FB} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h500} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b101, 12'h501} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b101, 12'h505} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h509} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'h50B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h50C} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b101, 12'h50D} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b101, 12'h50E} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h50F} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b101, 12'h510} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h511} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h513} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h514} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b101, 12'h515} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h516} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h517} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'h518} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h51C} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b101, 12'h51D} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h520} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h521} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b101, 12'h523} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h524} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b101, 12'h525} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h529} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b101, 12'h52B} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h52C} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h52D} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b101, 12'h52F} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h530} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b101, 12'h531} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h534} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b101, 12'h535} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h538} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b101, 12'h539} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h53C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b101, 12'h53D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h540} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b101, 12'h541} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h544} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b101, 12'h545} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h548} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b101, 12'h549} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h54C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b101, 12'h54D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h550} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b101, 12'h551} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h554} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b101, 12'h555} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h558} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b101, 12'h559} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h55C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b101, 12'h55D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h560} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b101, 12'h561} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h564} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b101, 12'h565} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h568} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b101, 12'h569} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h56C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b101, 12'h56D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h570} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b101, 12'h571} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h574} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b101, 12'h575} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h578} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b101, 12'h579} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h57C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b101, 12'h57D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h580} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b101, 12'h581} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h584} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b101, 12'h585} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h588} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b101, 12'h589} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h58C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b101, 12'h58D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h590} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b101, 12'h591} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h594} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b101, 12'h595} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h598} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b101, 12'h599} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h59C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b101, 12'h59D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b101, 12'h5A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b101, 12'h5A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b101, 12'h5A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b101, 12'h5AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b101, 12'h5B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b101, 12'h5B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b101, 12'h5B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b101, 12'h5BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5C0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b101, 12'h5C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b101, 12'h5C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5C8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b101, 12'h5C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5CC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b101, 12'h5CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5D0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b101, 12'h5D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5D4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b101, 12'h5D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5D8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b101, 12'h5D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b101, 12'h5DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b101, 12'h5E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b101, 12'h5E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5E8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b101, 12'h5E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5EC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b101, 12'h5ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b101, 12'h5F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5F4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b101, 12'h5F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5F8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b101, 12'h5F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h5FC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b101, 12'h5FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h600} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'h601} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h604} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b101, 12'h605} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h608} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'h609} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h60C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b101, 12'h60D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h610} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b101, 12'h611} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h614} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b101, 12'h615} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h618} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b101, 12'h619} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h61C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'h61D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h620} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b101, 12'h621} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h624} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b101, 12'h625} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h628} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b101, 12'h629} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h62C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b101, 12'h62D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h630} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b101, 12'h631} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h634} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b101, 12'h635} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h638} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b101, 12'h639} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h63C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b101, 12'h63D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h640} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'h641} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h644} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b101, 12'h645} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h648} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b101, 12'h649} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h64C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b101, 12'h64D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h650} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b101, 12'h651} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h654} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b101, 12'h655} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h658} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b101, 12'h659} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h65C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b101, 12'h65D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h660} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b101, 12'h661} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h664} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'h665} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h668} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b101, 12'h669} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h66C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b101, 12'h66D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h670} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b101, 12'h671} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h674} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b101, 12'h675} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h678} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b101, 12'h679} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h67C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b101, 12'h67D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h680} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'h681} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h684} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b101, 12'h685} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h688} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b101, 12'h689} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h68C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b101, 12'h68D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h690} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b101, 12'h691} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h694} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b101, 12'h695} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h698} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b101, 12'h699} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h69C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b101, 12'h69D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6A0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b101, 12'h6A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6A4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b101, 12'h6A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6A8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b101, 12'h6A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6AC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b101, 12'h6AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6B0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b101, 12'h6B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6B4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b101, 12'h6B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6B8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b101, 12'h6B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6BC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b101, 12'h6BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6C0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'h6C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6C4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b101, 12'h6C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6C8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b101, 12'h6C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6CC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b101, 12'h6CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6D0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b101, 12'h6D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6D4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b101, 12'h6D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6D8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b101, 12'h6D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6DC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b101, 12'h6DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6E0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b101, 12'h6E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6E4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b101, 12'h6E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6E8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b101, 12'h6E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6EC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b101, 12'h6ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6F0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b101, 12'h6F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6F4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b101, 12'h6F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6F8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b101, 12'h6F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h6FC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b101, 12'h6FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h700} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b101, 12'h701} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h704} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b101, 12'h705} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h708} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b101, 12'h709} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h70C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b101, 12'h70D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h710} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b101, 12'h711} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h714} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b101, 12'h715} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h718} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b101, 12'h719} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h71C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b101, 12'h71D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h720} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b101, 12'h721} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h724} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b101, 12'h725} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h728} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b101, 12'h729} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h72C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b101, 12'h72D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h730} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b101, 12'h731} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h734} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b101, 12'h735} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h738} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b101, 12'h739} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h73C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b101, 12'h73D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h740} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'h741} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h744} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b101, 12'h745} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h748} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b101, 12'h749} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h74C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b101, 12'h74D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h750} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b101, 12'h751} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h754} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b101, 12'h755} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h758} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b101, 12'h759} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h75C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b101, 12'h75D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h760} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b101, 12'h761} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h764} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b101, 12'h765} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h768} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b101, 12'h769} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h76C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b101, 12'h76D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h770} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b101, 12'h771} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h774} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b101, 12'h775} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h778} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b101, 12'h779} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h77C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b101, 12'h77D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h780} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'h781} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h784} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b101, 12'h785} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h788} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b101, 12'h789} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h78C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b101, 12'h78D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h790} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b101, 12'h791} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h794} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b101, 12'h795} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h798} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b101, 12'h799} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h79C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b101, 12'h79D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7A0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'h7A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7A4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b101, 12'h7A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7A8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b101, 12'h7A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7AC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b101, 12'h7AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7B0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b101, 12'h7B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7B4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b101, 12'h7B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7B8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b101, 12'h7B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7BC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b101, 12'h7BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7C0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b101, 12'h7C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7C4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b101, 12'h7C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7C8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b101, 12'h7C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7CC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b101, 12'h7CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7D0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b101, 12'h7D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7D4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b101, 12'h7D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7D8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b101, 12'h7D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7DC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b101, 12'h7DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7E0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b101, 12'h7E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7E4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b101, 12'h7E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7E8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b101, 12'h7E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7EC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b101, 12'h7ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7F0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b101, 12'h7F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7F4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b101, 12'h7F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7F8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b101, 12'h7F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h7FC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b101, 12'h7FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h801} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h804} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'h805} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h808} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'h809} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h80C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'h80D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h810} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'h811} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h814} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b101, 12'h815} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h818} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b101, 12'h819} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h81C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'h81D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h820} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b101, 12'h821} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h824} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'h825} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h828} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b101, 12'h829} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h82C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'h82D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h830} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b101, 12'h831} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h834} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b101, 12'h835} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h838} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'h839} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h83C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'h83D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h840} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h841} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h844} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b101, 12'h845} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h848} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b101, 12'h849} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h84C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b101, 12'h84D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h850} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b101, 12'h851} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h854} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b101, 12'h855} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h858} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b101, 12'h859} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h85C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b101, 12'h85D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h860} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b101, 12'h861} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h864} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b101, 12'h865} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h868} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b101, 12'h869} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h86C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b101, 12'h86D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h870} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b101, 12'h871} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h874} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b101, 12'h875} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h878} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b101, 12'h879} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h87C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'h87D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h880} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'h881} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h884} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b101, 12'h885} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h888} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'h889} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h88C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b101, 12'h88D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h890} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b101, 12'h891} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h894} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b101, 12'h895} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h898} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b101, 12'h899} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h89C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b101, 12'h89D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8A0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b101, 12'h8A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8A4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'h8A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8A8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b101, 12'h8A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8AC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b101, 12'h8AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8B0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'h8B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8B4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b101, 12'h8B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8B8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b101, 12'h8B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8BC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'h8BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8C0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b101, 12'h8C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8C4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b101, 12'h8C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8C8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b101, 12'h8C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8CC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b101, 12'h8CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8D0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b101, 12'h8D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8D4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b101, 12'h8D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8D8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b101, 12'h8D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8DC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b101, 12'h8DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8E0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b101, 12'h8E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8E4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b101, 12'h8E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8E8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b101, 12'h8E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8EC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b101, 12'h8ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8F0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b101, 12'h8F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8F4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b101, 12'h8F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b101, 12'h8F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h8FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b101, 12'h8FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h900} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'h901} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h904} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b101, 12'h905} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h908} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b101, 12'h909} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h90C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b101, 12'h90D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h910} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b101, 12'h911} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h914} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b101, 12'h915} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h918} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b101, 12'h919} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h91C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b101, 12'h91D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h920} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b101, 12'h921} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h924} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b101, 12'h925} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h928} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b101, 12'h929} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h92C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b101, 12'h92D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h930} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b101, 12'h931} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h934} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b101, 12'h935} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h938} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b101, 12'h939} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h93C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b101, 12'h93D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h940} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b101, 12'h941} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h944} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b101, 12'h945} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h948} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b101, 12'h949} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h94C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b101, 12'h94D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h950} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b101, 12'h951} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h954} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b101, 12'h955} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h958} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b101, 12'h959} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h95C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b101, 12'h95D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h960} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b101, 12'h961} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h964} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b101, 12'h965} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h968} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b101, 12'h969} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h96C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b101, 12'h96D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h970} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b101, 12'h971} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h974} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b101, 12'h975} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h978} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b101, 12'h979} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h97C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b101, 12'h97D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h980} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b101, 12'h981} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h984} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b101, 12'h985} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h988} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b101, 12'h989} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h98C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b101, 12'h98D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h990} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b101, 12'h991} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h994} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b101, 12'h995} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h998} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b101, 12'h999} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h99C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b101, 12'h99D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b101, 12'h9A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b101, 12'h9A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b101, 12'h9A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b101, 12'h9AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b101, 12'h9B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b101, 12'h9B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b101, 12'h9B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b101, 12'h9BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9C0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b101, 12'h9C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b101, 12'h9C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9C8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b101, 12'h9C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9CC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b101, 12'h9CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9D0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b101, 12'h9D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9D4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b101, 12'h9D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9D8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b101, 12'h9D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b101, 12'h9DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b101, 12'h9E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b101, 12'h9E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9E8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b101, 12'h9E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9EC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b101, 12'h9ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b101, 12'h9F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9F4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b101, 12'h9F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9F8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b101, 12'h9F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'h9FC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b101, 12'h9FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA00} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'hA01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA04} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b101, 12'hA05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA08} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'hA09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA0C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b101, 12'hA0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA10} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b101, 12'hA11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA14} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b101, 12'hA15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA18} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b101, 12'hA19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA1C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'hA1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA20} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b101, 12'hA21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA24} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b101, 12'hA25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA28} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b101, 12'hA29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA2C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b101, 12'hA2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA30} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b101, 12'hA31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA34} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b101, 12'hA35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA38} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b101, 12'hA39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA3C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b101, 12'hA3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA40} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'hA41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA44} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b101, 12'hA45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA48} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b101, 12'hA49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA4C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b101, 12'hA4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA50} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b101, 12'hA51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA54} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b101, 12'hA55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA58} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b101, 12'hA59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA5C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b101, 12'hA5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA60} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b101, 12'hA61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA64} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'hA65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA68} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b101, 12'hA69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA6C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b101, 12'hA6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA70} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b101, 12'hA71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA74} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b101, 12'hA75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b101, 12'hA79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA7C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b101, 12'hA7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA80} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'hA81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA84} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b101, 12'hA85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA88} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b101, 12'hA89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA8C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b101, 12'hA8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA90} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b101, 12'hA91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA94} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b101, 12'hA95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA98} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b101, 12'hA99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hA9C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b101, 12'hA9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAA0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b101, 12'hAA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAA4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b101, 12'hAA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAA8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b101, 12'hAA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAAC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b101, 12'hAAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAB0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b101, 12'hAB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAB4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b101, 12'hAB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAB8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b101, 12'hAB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hABC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b101, 12'hABD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAC0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'hAC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAC4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b101, 12'hAC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAC8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b101, 12'hAC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hACC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b101, 12'hACD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAD0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b101, 12'hAD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAD4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b101, 12'hAD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAD8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b101, 12'hAD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hADC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b101, 12'hADD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAE0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b101, 12'hAE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAE4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b101, 12'hAE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAE8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b101, 12'hAE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAEC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b101, 12'hAED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAF0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b101, 12'hAF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAF4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b101, 12'hAF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAF8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b101, 12'hAF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hAFC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b101, 12'hAFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB00} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b101, 12'hB01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB04} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b101, 12'hB05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB08} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b101, 12'hB09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB0C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b101, 12'hB0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB10} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b101, 12'hB11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB14} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b101, 12'hB15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB18} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b101, 12'hB19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB1C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b101, 12'hB1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB20} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b101, 12'hB21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB24} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b101, 12'hB25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB28} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b101, 12'hB29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB2C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b101, 12'hB2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB30} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b101, 12'hB31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB34} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b101, 12'hB35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB38} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b101, 12'hB39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB3C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b101, 12'hB3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB40} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'hB41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB44} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b101, 12'hB45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB48} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b101, 12'hB49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB4C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b101, 12'hB4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB50} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b101, 12'hB51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB54} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b101, 12'hB55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB58} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b101, 12'hB59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB5C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b101, 12'hB5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB60} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b101, 12'hB61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB64} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b101, 12'hB65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB68} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b101, 12'hB69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB6C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b101, 12'hB6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB70} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b101, 12'hB71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB74} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b101, 12'hB75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB78} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b101, 12'hB79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB7C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b101, 12'hB7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB80} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'hB81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB84} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b101, 12'hB85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB88} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b101, 12'hB89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB8C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b101, 12'hB8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB90} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b101, 12'hB91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB94} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b101, 12'hB95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB98} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b101, 12'hB99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hB9C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b101, 12'hB9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBA0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'hBA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBA4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b101, 12'hBA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBA8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b101, 12'hBA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBAC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b101, 12'hBAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBB0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b101, 12'hBB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBB4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b101, 12'hBB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBB8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b101, 12'hBB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBBC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b101, 12'hBBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBC0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b101, 12'hBC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBC4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b101, 12'hBC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBC8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b101, 12'hBC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBCC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b101, 12'hBCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBD0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b101, 12'hBD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBD4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b101, 12'hBD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBD8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b101, 12'hBD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBDC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b101, 12'hBDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBE0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b101, 12'hBE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBE4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b101, 12'hBE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBE8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b101, 12'hBE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBEC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b101, 12'hBED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBF0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b101, 12'hBF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBF4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b101, 12'hBF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBF8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b101, 12'hBF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hBFC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b101, 12'hBFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC04} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b101, 12'hC05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC08} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b101, 12'hC09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC0C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b101, 12'hC0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC10} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b101, 12'hC11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC14} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b101, 12'hC15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC18} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b101, 12'hC19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC1C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b101, 12'hC1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC20} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b101, 12'hC21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC24} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b101, 12'hC25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC28} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b101, 12'hC29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC2C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b101, 12'hC2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC30} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b101, 12'hC31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC34} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b101, 12'hC35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC38} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b101, 12'hC39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC3C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b101, 12'hC3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC40} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC44} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b101, 12'hC45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC48} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b101, 12'hC49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC4C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b101, 12'hC4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC50} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b101, 12'hC51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC54} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b101, 12'hC55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC58} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b101, 12'hC59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC5C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b101, 12'hC5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC60} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b101, 12'hC61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC64} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b101, 12'hC65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC68} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b101, 12'hC69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC6C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b101, 12'hC6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC70} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b101, 12'hC71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC74} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b101, 12'hC75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC78} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b101, 12'hC79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC7C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b101, 12'hC7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC80} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b101, 12'hC81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC84} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b101, 12'hC85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC88} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b101, 12'hC89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC8C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b101, 12'hC8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC90} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b101, 12'hC91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC94} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b101, 12'hC95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC98} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b101, 12'hC99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hC9C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b101, 12'hC9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCA0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b101, 12'hCA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCA4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b101, 12'hCA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCA8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b101, 12'hCA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCAC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b101, 12'hCAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCB0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b101, 12'hCB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCB4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b101, 12'hCB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCB8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b101, 12'hCB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCBC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b101, 12'hCBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCC0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b101, 12'hCC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCC4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b101, 12'hCC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCC8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b101, 12'hCC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCCC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b101, 12'hCCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCD0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b101, 12'hCD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCD4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b101, 12'hCD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCD8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b101, 12'hCD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCDC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b101, 12'hCDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCE0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b101, 12'hCE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCE4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b101, 12'hCE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCE8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b101, 12'hCE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCEC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b101, 12'hCED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCF0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b101, 12'hCF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCF4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b101, 12'hCF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCF8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b101, 12'hCF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hCFC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b101, 12'hCFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD00} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b101, 12'hD01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD04} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b101, 12'hD05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD08} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b101, 12'hD09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD0C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b101, 12'hD0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD10} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b101, 12'hD11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD14} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b101, 12'hD15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD18} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b101, 12'hD19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD1C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b101, 12'hD1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD20} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b101, 12'hD21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD24} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b101, 12'hD25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD28} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b101, 12'hD29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD2C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b101, 12'hD2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD30} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b101, 12'hD31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD34} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b101, 12'hD35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD38} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b101, 12'hD39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD3C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b101, 12'hD3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD40} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b101, 12'hD41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD44} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b101, 12'hD45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD48} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b101, 12'hD49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD4C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b101, 12'hD4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD50} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b101, 12'hD51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD54} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b101, 12'hD55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD58} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b101, 12'hD59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD5C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b101, 12'hD5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD60} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b101, 12'hD61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD64} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b101, 12'hD65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD68} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b101, 12'hD69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD6C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b101, 12'hD6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD70} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b101, 12'hD71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD74} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b101, 12'hD75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD78} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b101, 12'hD79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD7C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b101, 12'hD7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD80} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b101, 12'hD81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD84} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b101, 12'hD85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD88} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b101, 12'hD89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD8C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b101, 12'hD8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD90} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b101, 12'hD91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD94} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b101, 12'hD95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD98} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b101, 12'hD99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hD9C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b101, 12'hD9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDA0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b101, 12'hDA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDA4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b101, 12'hDA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDA8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b101, 12'hDA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDAC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b101, 12'hDAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDB0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b101, 12'hDB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDB4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b101, 12'hDB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDB8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b101, 12'hDB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDBC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b101, 12'hDBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDC0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b101, 12'hDC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDC4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b101, 12'hDC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDC8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b101, 12'hDC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDCC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b101, 12'hDCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDD0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b101, 12'hDD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDD4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b101, 12'hDD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDD8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b101, 12'hDD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDDC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b101, 12'hDDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDE0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b101, 12'hDE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDE4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b101, 12'hDE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDE8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b101, 12'hDE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDEC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b101, 12'hDED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDF0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b101, 12'hDF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDF4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b101, 12'hDF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDF8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b101, 12'hDF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hDFC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b101, 12'hDFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE00} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b101, 12'hE01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE04} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b101, 12'hE05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE08} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b101, 12'hE09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE0C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b101, 12'hE0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE10} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b101, 12'hE11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE14} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b101, 12'hE15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE18} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b101, 12'hE19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE1C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b101, 12'hE1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE20} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b101, 12'hE21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE24} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b101, 12'hE25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE28} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b101, 12'hE29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE2C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b101, 12'hE2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE30} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b101, 12'hE31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE34} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b101, 12'hE35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE38} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b101, 12'hE39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE3C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b101, 12'hE3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE40} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b101, 12'hE41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE44} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b101, 12'hE45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE48} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b101, 12'hE49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE4C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b101, 12'hE4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE50} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b101, 12'hE51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE54} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b101, 12'hE55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE58} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b101, 12'hE59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE5C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b101, 12'hE5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE60} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b101, 12'hE61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE64} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b101, 12'hE65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE68} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b101, 12'hE69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE6C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b101, 12'hE6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE70} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b101, 12'hE71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE74} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b101, 12'hE75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b101, 12'hE79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE7C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b101, 12'hE7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE80} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b101, 12'hE81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE84} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b101, 12'hE85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE88} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b101, 12'hE89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE8C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b101, 12'hE8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE90} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b101, 12'hE91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE94} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b101, 12'hE95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE98} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b101, 12'hE99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hE9C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b101, 12'hE9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEA0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b101, 12'hEA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEA4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b101, 12'hEA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEA8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b101, 12'hEA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEAC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b101, 12'hEAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEB0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b101, 12'hEB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEB4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b101, 12'hEB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEB8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b101, 12'hEB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEBC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b101, 12'hEBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEC0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b101, 12'hEC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEC4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b101, 12'hEC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEC8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b101, 12'hEC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hECC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b101, 12'hECD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hED0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b101, 12'hED1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hED4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b101, 12'hED5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hED8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b101, 12'hED9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEDC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b101, 12'hEDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEE0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b101, 12'hEE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEE4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b101, 12'hEE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEE8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b101, 12'hEE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEEC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b101, 12'hEED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEF0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b101, 12'hEF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEF4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b101, 12'hEF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEF8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b101, 12'hEF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hEFC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b101, 12'hEFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF00} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b101, 12'hF01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF04} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b101, 12'hF05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF08} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b101, 12'hF09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF0C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b101, 12'hF0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF10} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b101, 12'hF11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF14} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b101, 12'hF15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF18} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b101, 12'hF19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF1C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b101, 12'hF1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF20} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b101, 12'hF21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF24} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b101, 12'hF25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF28} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b101, 12'hF29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF2C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b101, 12'hF2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF30} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b101, 12'hF31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF34} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b101, 12'hF35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF38} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b101, 12'hF39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF3C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b101, 12'hF3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF40} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b101, 12'hF41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF44} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b101, 12'hF45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF48} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b101, 12'hF49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF4C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b101, 12'hF4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF50} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b101, 12'hF51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF54} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b101, 12'hF55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF58} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b101, 12'hF59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF5C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b101, 12'hF5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF60} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b101, 12'hF61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF64} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b101, 12'hF65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF68} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b101, 12'hF69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF6C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b101, 12'hF6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF70} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b101, 12'hF71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF74} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b101, 12'hF75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF78} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b101, 12'hF79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF7C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b101, 12'hF7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF80} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b101, 12'hF81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF84} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b101, 12'hF85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF88} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b101, 12'hF89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF8C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b101, 12'hF8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF90} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b101, 12'hF91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF94} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b101, 12'hF95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF98} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b101, 12'hF99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hF9C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b101, 12'hF9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFA0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b101, 12'hFA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFA4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b101, 12'hFA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFA8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b101, 12'hFA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFAC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b101, 12'hFAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFB0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b101, 12'hFB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFB4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b101, 12'hFB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFB8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b101, 12'hFB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFBC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b101, 12'hFBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFC0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b101, 12'hFC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFC4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b101, 12'hFC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFC8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b101, 12'hFC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFCC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b101, 12'hFCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFD0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b101, 12'hFD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFD4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b101, 12'hFD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFD8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b101, 12'hFD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFDC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b101, 12'hFDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFE0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b101, 12'hFE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFE4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b101, 12'hFE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFE8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b101, 12'hFE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFEC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b101, 12'hFED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFF0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b101, 12'hFF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFF4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b101, 12'hFF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFF8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b101, 12'hFF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b101, 12'hFFC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b101, 12'hFFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h001} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h004} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b110, 12'h005} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h008} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b110, 12'h009} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h00C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b110, 12'h00D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h010} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b110, 12'h011} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h014} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b110, 12'h015} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h018} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b110, 12'h019} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h01C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b110, 12'h01D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h020} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b110, 12'h021} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h024} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b110, 12'h025} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h028} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b110, 12'h029} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h02C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b110, 12'h02D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h030} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b110, 12'h031} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h034} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b110, 12'h035} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h038} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b110, 12'h039} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h03C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b110, 12'h03D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h040} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h041} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h044} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b110, 12'h045} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h048} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b110, 12'h049} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h04C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b110, 12'h04D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h050} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b110, 12'h051} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h054} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b110, 12'h055} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h058} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b110, 12'h059} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h05C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b110, 12'h05D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h060} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b110, 12'h061} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h064} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b110, 12'h065} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h068} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b110, 12'h069} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h06C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b110, 12'h06D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h070} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b110, 12'h071} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h074} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b110, 12'h075} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h078} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b110, 12'h079} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h07C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b110, 12'h07D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h080} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b110, 12'h081} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h084} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b110, 12'h085} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h088} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b110, 12'h089} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h08C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b110, 12'h08D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h090} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b110, 12'h091} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h094} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b110, 12'h095} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h098} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b110, 12'h099} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h09C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b110, 12'h09D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0A0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b110, 12'h0A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0A4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b110, 12'h0A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0A8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b110, 12'h0A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0AC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b110, 12'h0AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0B0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b110, 12'h0B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0B4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b110, 12'h0B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0B8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b110, 12'h0B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0BC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b110, 12'h0BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0C0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b110, 12'h0C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0C4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b110, 12'h0C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0C8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b110, 12'h0C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0CC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b110, 12'h0CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0D0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b110, 12'h0D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0D4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b110, 12'h0D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0D8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b110, 12'h0D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0DC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b110, 12'h0DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0E0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b110, 12'h0E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0E4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b110, 12'h0E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0E8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b110, 12'h0E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0EC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b110, 12'h0ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0F0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b110, 12'h0F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0F4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b110, 12'h0F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b110, 12'h0F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h0FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b110, 12'h0FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h100} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b110, 12'h101} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h104} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b110, 12'h105} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h108} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b110, 12'h109} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h10C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b110, 12'h10D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h110} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b110, 12'h111} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h114} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b110, 12'h115} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h118} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b110, 12'h119} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h11C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b110, 12'h11D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h120} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b110, 12'h121} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h124} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b110, 12'h125} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h128} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b110, 12'h129} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h12C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b110, 12'h12D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h130} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b110, 12'h131} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h134} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b110, 12'h135} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h138} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b110, 12'h139} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h13C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b110, 12'h13D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h140} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b110, 12'h141} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h144} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b110, 12'h145} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h148} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b110, 12'h149} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h14C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b110, 12'h14D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h150} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b110, 12'h151} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h154} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b110, 12'h155} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h158} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b110, 12'h159} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h15C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b110, 12'h15D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h160} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b110, 12'h161} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h164} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b110, 12'h165} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h168} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b110, 12'h169} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h16C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b110, 12'h16D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h170} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b110, 12'h171} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h174} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b110, 12'h175} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h178} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b110, 12'h179} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h17C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b110, 12'h17D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h180} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b110, 12'h181} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h184} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b110, 12'h185} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h188} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b110, 12'h189} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h18C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b110, 12'h18D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h190} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b110, 12'h191} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h194} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b110, 12'h195} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h198} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b110, 12'h199} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h19C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b110, 12'h19D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b110, 12'h1A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b110, 12'h1A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b110, 12'h1A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b110, 12'h1AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b110, 12'h1B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b110, 12'h1B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b110, 12'h1B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b110, 12'h1BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1C0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b110, 12'h1C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b110, 12'h1C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1C8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b110, 12'h1C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1CC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b110, 12'h1CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1D0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b110, 12'h1D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1D4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b110, 12'h1D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1D8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b110, 12'h1D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b110, 12'h1DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b110, 12'h1E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b110, 12'h1E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1E8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b110, 12'h1E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1EC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b110, 12'h1ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b110, 12'h1F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1F4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b110, 12'h1F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1F8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b110, 12'h1F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h1FC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b110, 12'h1FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h200} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b110, 12'h201} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h204} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b110, 12'h205} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h208} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b110, 12'h209} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h20C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b110, 12'h20D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h210} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b110, 12'h211} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h214} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b110, 12'h215} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h218} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b110, 12'h219} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h21C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b110, 12'h21D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h220} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b110, 12'h221} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h224} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b110, 12'h225} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h228} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b110, 12'h229} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h22C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b110, 12'h22D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h230} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b110, 12'h231} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h234} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b110, 12'h235} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h238} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b110, 12'h239} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h23C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b110, 12'h23D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h240} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b110, 12'h241} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h244} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b110, 12'h245} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h248} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b110, 12'h249} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h24C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b110, 12'h24D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h250} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b110, 12'h251} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h254} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b110, 12'h255} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h258} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b110, 12'h259} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h25C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b110, 12'h25D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h260} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b110, 12'h261} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h264} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b110, 12'h265} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h268} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b110, 12'h269} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h26C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b110, 12'h26D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h270} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b110, 12'h271} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h274} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b110, 12'h275} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h278} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b110, 12'h279} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h27C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b110, 12'h27D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h280} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b110, 12'h281} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h284} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b110, 12'h285} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h288} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b110, 12'h289} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h28C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b110, 12'h28D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h290} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b110, 12'h291} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h294} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b110, 12'h295} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h298} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b110, 12'h299} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h29C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b110, 12'h29D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2A0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b110, 12'h2A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2A4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b110, 12'h2A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2A8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b110, 12'h2A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2AC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b110, 12'h2AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2B0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b110, 12'h2B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2B4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b110, 12'h2B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2B8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b110, 12'h2B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2BC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b110, 12'h2BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2C0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b110, 12'h2C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2C4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b110, 12'h2C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2C8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b110, 12'h2C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2CC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b110, 12'h2CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2D0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b110, 12'h2D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2D4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b110, 12'h2D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2D8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b110, 12'h2D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2DC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b110, 12'h2DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2E0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b110, 12'h2E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2E4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b110, 12'h2E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2E8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b110, 12'h2E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2EC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b110, 12'h2ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2F0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b110, 12'h2F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2F4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b110, 12'h2F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2F8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b110, 12'h2F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h2FC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b110, 12'h2FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h300} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b110, 12'h301} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h304} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b110, 12'h305} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h308} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b110, 12'h309} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h30C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b110, 12'h30D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h310} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b110, 12'h311} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h314} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b110, 12'h315} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h318} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b110, 12'h319} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h31C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b110, 12'h31D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h320} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b110, 12'h321} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h324} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b110, 12'h325} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h328} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b110, 12'h329} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h32C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b110, 12'h32D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h330} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b110, 12'h331} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h334} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b110, 12'h335} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h338} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b110, 12'h339} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h33C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b110, 12'h33D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h340} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b110, 12'h341} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h344} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b110, 12'h345} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h348} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b110, 12'h349} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h34C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b110, 12'h34D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h350} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b110, 12'h351} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h354} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b110, 12'h355} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h358} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b110, 12'h359} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h35C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b110, 12'h35D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h360} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b110, 12'h361} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h364} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b110, 12'h365} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h368} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b110, 12'h369} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h36C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b110, 12'h36D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h370} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b110, 12'h371} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h374} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b110, 12'h375} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h378} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b110, 12'h379} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h37C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b110, 12'h37D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h380} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b110, 12'h381} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h384} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b110, 12'h385} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h388} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b110, 12'h389} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h38C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b110, 12'h38D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h390} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b110, 12'h391} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h394} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b110, 12'h395} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h398} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b110, 12'h399} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h39C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b110, 12'h39D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3A0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b110, 12'h3A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3A4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b110, 12'h3A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3A8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b110, 12'h3A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3AC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b110, 12'h3AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3B0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b110, 12'h3B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3B4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b110, 12'h3B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3B8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b110, 12'h3B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3BC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b110, 12'h3BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3C0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b110, 12'h3C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3C4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b110, 12'h3C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3C8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b110, 12'h3C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3CC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b110, 12'h3CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3D0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b110, 12'h3D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3D4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b110, 12'h3D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3D8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b110, 12'h3D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3DC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b110, 12'h3DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3E0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b110, 12'h3E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3E4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b110, 12'h3E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3E8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b110, 12'h3E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3EC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b110, 12'h3ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3F0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b110, 12'h3F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3F4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b110, 12'h3F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3F8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b110, 12'h3F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h3FC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b110, 12'h3FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h401} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h404} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b110, 12'h405} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h408} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b110, 12'h409} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h40C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b110, 12'h40D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h410} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b110, 12'h411} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h414} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b110, 12'h415} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h418} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b110, 12'h419} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h41C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b110, 12'h41D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h420} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b110, 12'h421} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h424} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b110, 12'h425} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h428} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b110, 12'h429} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h42C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b110, 12'h42D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h430} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b110, 12'h431} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h434} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b110, 12'h435} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h438} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b110, 12'h439} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h43C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b110, 12'h43D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h440} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h441} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h444} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b110, 12'h445} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h448} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b110, 12'h449} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h44C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b110, 12'h44D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h450} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b110, 12'h451} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h454} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b110, 12'h455} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h458} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b110, 12'h459} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h45C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b110, 12'h45D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h460} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b110, 12'h461} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h464} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b110, 12'h465} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h468} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b110, 12'h469} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h46C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b110, 12'h46D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h470} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b110, 12'h471} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h474} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b110, 12'h475} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h478} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b110, 12'h479} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h47C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b110, 12'h47D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h480} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b110, 12'h481} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h484} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b110, 12'h485} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h488} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b110, 12'h489} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h48C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b110, 12'h48D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h490} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b110, 12'h491} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h494} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b110, 12'h495} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h498} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b110, 12'h499} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h49C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b110, 12'h49D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4A0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b110, 12'h4A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4A4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b110, 12'h4A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4A8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b110, 12'h4A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4AC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b110, 12'h4AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4B0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b110, 12'h4B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4B4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b110, 12'h4B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4B8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b110, 12'h4B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4BC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b110, 12'h4BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4C0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b110, 12'h4C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4C4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b110, 12'h4C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4C8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b110, 12'h4C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4CC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b110, 12'h4CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4D0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b110, 12'h4D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4D4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b110, 12'h4D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4D8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b110, 12'h4D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4DC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b110, 12'h4DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4E0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b110, 12'h4E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4E4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b110, 12'h4E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4E8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b110, 12'h4E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4EC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b110, 12'h4ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4F0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b110, 12'h4F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4F4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b110, 12'h4F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b110, 12'h4F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h4FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b110, 12'h4FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h500} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b110, 12'h501} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h504} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b110, 12'h505} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h508} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b110, 12'h509} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h50C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b110, 12'h50D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h510} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b110, 12'h511} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h514} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b110, 12'h515} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h518} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b110, 12'h519} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h51C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b110, 12'h51D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h520} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b110, 12'h521} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h524} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b110, 12'h525} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h528} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b110, 12'h529} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h52C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b110, 12'h52D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h530} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b110, 12'h531} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h534} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b110, 12'h535} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h538} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b110, 12'h539} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h53C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b110, 12'h53D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h540} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b110, 12'h541} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h544} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b110, 12'h545} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h548} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b110, 12'h549} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h54C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b110, 12'h54D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h550} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b110, 12'h551} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h554} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b110, 12'h555} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h558} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b110, 12'h559} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h55C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b110, 12'h55D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h560} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b110, 12'h561} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h564} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b110, 12'h565} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h568} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b110, 12'h569} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h56C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b110, 12'h56D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h570} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b110, 12'h571} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h574} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b110, 12'h575} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h578} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b110, 12'h579} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h57C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b110, 12'h57D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h580} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b110, 12'h581} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h584} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b110, 12'h585} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h588} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b110, 12'h589} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h58C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b110, 12'h58D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h590} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b110, 12'h591} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h594} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b110, 12'h595} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h598} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b110, 12'h599} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h59C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b110, 12'h59D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b110, 12'h5A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b110, 12'h5A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b110, 12'h5A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b110, 12'h5AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b110, 12'h5B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b110, 12'h5B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b110, 12'h5B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b110, 12'h5BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5C0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b110, 12'h5C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b110, 12'h5C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5C8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b110, 12'h5C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5CC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b110, 12'h5CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5D0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b110, 12'h5D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5D4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b110, 12'h5D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5D8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b110, 12'h5D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b110, 12'h5DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b110, 12'h5E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b110, 12'h5E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5E8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b110, 12'h5E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5EC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b110, 12'h5ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b110, 12'h5F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5F4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b110, 12'h5F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5F8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b110, 12'h5F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h5FC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b110, 12'h5FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h600} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b110, 12'h601} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h604} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b110, 12'h605} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h608} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b110, 12'h609} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h60C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b110, 12'h60D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h610} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b110, 12'h611} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h614} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b110, 12'h615} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h618} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b110, 12'h619} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h61C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b110, 12'h61D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h620} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b110, 12'h621} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h624} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b110, 12'h625} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h628} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b110, 12'h629} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h62C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b110, 12'h62D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h630} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b110, 12'h631} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h634} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b110, 12'h635} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h638} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b110, 12'h639} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h63C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b110, 12'h63D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h640} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b110, 12'h641} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h644} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b110, 12'h645} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h648} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b110, 12'h649} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h64C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b110, 12'h64D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h650} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b110, 12'h651} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h654} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b110, 12'h655} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h658} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b110, 12'h659} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h65C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b110, 12'h65D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h660} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b110, 12'h661} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h664} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b110, 12'h665} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h668} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b110, 12'h669} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h66C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b110, 12'h66D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h670} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b110, 12'h671} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h674} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b110, 12'h675} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h678} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b110, 12'h679} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h67C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b110, 12'h67D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h680} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b110, 12'h681} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h684} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b110, 12'h685} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h688} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b110, 12'h689} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h68C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b110, 12'h68D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h690} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b110, 12'h691} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h694} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b110, 12'h695} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h698} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b110, 12'h699} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h69C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b110, 12'h69D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6A0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b110, 12'h6A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6A4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b110, 12'h6A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6A8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b110, 12'h6A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6AC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b110, 12'h6AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6B0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b110, 12'h6B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6B4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b110, 12'h6B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6B8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b110, 12'h6B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6BC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b110, 12'h6BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6C0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b110, 12'h6C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6C4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b110, 12'h6C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6C8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b110, 12'h6C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6CC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b110, 12'h6CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6D0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b110, 12'h6D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6D4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b110, 12'h6D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6D8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b110, 12'h6D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6DC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b110, 12'h6DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6E0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b110, 12'h6E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6E4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b110, 12'h6E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6E8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b110, 12'h6E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6EC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b110, 12'h6ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6F0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b110, 12'h6F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6F4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b110, 12'h6F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6F8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b110, 12'h6F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h6FC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b110, 12'h6FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h700} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b110, 12'h701} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h704} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b110, 12'h705} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h708} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b110, 12'h709} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h70C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b110, 12'h70D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h710} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b110, 12'h711} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h714} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b110, 12'h715} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h718} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b110, 12'h719} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h71C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b110, 12'h71D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h720} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b110, 12'h721} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h724} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b110, 12'h725} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h728} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b110, 12'h729} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h72C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b110, 12'h72D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h730} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b110, 12'h731} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h734} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b110, 12'h735} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h738} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b110, 12'h739} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h73C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b110, 12'h73D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h740} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b110, 12'h741} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h744} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b110, 12'h745} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h748} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b110, 12'h749} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h74C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b110, 12'h74D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h750} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b110, 12'h751} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h754} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b110, 12'h755} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h758} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b110, 12'h759} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h75C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b110, 12'h75D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h760} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b110, 12'h761} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h764} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b110, 12'h765} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h768} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b110, 12'h769} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h76C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b110, 12'h76D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h770} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b110, 12'h771} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h774} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b110, 12'h775} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h778} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b110, 12'h779} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h77C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b110, 12'h77D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h780} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b110, 12'h781} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h784} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b110, 12'h785} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h788} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b110, 12'h789} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h78C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b110, 12'h78D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h790} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b110, 12'h791} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h794} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b110, 12'h795} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h798} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b110, 12'h799} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h79C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b110, 12'h79D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7A0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b110, 12'h7A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7A4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b110, 12'h7A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7A8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b110, 12'h7A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7AC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b110, 12'h7AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7B0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b110, 12'h7B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7B4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b110, 12'h7B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7B8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b110, 12'h7B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7BC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b110, 12'h7BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7C0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b110, 12'h7C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7C4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b110, 12'h7C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7C8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b110, 12'h7C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7CC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b110, 12'h7CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7D0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b110, 12'h7D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7D4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b110, 12'h7D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7D8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b110, 12'h7D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7DC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b110, 12'h7DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7E0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b110, 12'h7E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7E4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b110, 12'h7E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7E8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b110, 12'h7E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7EC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b110, 12'h7ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7F0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b110, 12'h7F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7F4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b110, 12'h7F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7F8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b110, 12'h7F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h7FC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b110, 12'h7FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h801} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h804} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b110, 12'h805} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h808} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b110, 12'h809} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h80C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b110, 12'h80D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h810} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b110, 12'h811} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h814} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b110, 12'h815} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h818} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b110, 12'h819} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h81C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b110, 12'h81D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h820} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b110, 12'h821} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h824} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b110, 12'h825} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h828} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b110, 12'h829} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h82C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b110, 12'h82D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h830} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b110, 12'h831} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h834} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b110, 12'h835} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h838} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b110, 12'h839} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h83C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b110, 12'h83D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h840} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h841} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h844} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b110, 12'h845} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h848} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b110, 12'h849} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h84C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b110, 12'h84D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h850} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b110, 12'h851} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h854} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b110, 12'h855} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h858} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b110, 12'h859} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h85C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b110, 12'h85D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h860} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b110, 12'h861} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h864} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b110, 12'h865} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h868} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b110, 12'h869} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h86C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b110, 12'h86D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h870} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b110, 12'h871} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h874} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b110, 12'h875} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h878} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b110, 12'h879} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h87C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b110, 12'h87D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h880} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b110, 12'h881} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h884} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b110, 12'h885} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h888} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b110, 12'h889} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h88C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b110, 12'h88D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h890} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b110, 12'h891} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h894} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b110, 12'h895} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h898} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b110, 12'h899} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h89C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b110, 12'h89D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8A0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b110, 12'h8A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8A4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b110, 12'h8A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8A8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b110, 12'h8A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8AC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b110, 12'h8AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8B0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b110, 12'h8B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8B4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b110, 12'h8B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8B8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b110, 12'h8B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8BC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b110, 12'h8BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8C0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b110, 12'h8C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8C4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b110, 12'h8C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8C8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b110, 12'h8C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8CC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b110, 12'h8CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8D0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b110, 12'h8D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8D4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b110, 12'h8D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8D8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b110, 12'h8D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8DC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b110, 12'h8DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8E0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b110, 12'h8E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8E4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b110, 12'h8E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8E8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b110, 12'h8E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8EC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b110, 12'h8ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8F0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b110, 12'h8F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8F4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b110, 12'h8F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b110, 12'h8F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h8FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b110, 12'h8FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h900} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b110, 12'h901} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h904} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b110, 12'h905} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h908} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b110, 12'h909} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h90C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b110, 12'h90D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h910} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b110, 12'h911} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h914} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b110, 12'h915} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h918} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b110, 12'h919} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h91C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b110, 12'h91D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h920} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b110, 12'h921} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h924} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b110, 12'h925} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h928} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b110, 12'h929} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h92C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b110, 12'h92D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h930} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b110, 12'h931} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h934} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b110, 12'h935} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h938} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b110, 12'h939} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h93C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b110, 12'h93D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h940} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b110, 12'h941} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h944} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b110, 12'h945} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h948} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b110, 12'h949} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h94C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b110, 12'h94D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h950} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b110, 12'h951} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h954} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b110, 12'h955} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h958} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b110, 12'h959} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h95C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b110, 12'h95D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h960} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b110, 12'h961} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h964} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b110, 12'h965} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h968} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b110, 12'h969} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h96C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b110, 12'h96D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h970} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b110, 12'h971} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h974} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b110, 12'h975} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h978} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b110, 12'h979} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h97C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b110, 12'h97D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h980} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b110, 12'h981} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h984} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b110, 12'h985} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h988} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b110, 12'h989} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h98C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b110, 12'h98D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h990} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b110, 12'h991} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h994} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b110, 12'h995} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h998} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b110, 12'h999} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h99C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b110, 12'h99D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b110, 12'h9A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b110, 12'h9A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b110, 12'h9A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b110, 12'h9AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b110, 12'h9B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b110, 12'h9B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b110, 12'h9B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b110, 12'h9BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9C0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b110, 12'h9C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b110, 12'h9C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9C8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b110, 12'h9C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9CC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b110, 12'h9CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9D0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b110, 12'h9D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9D4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b110, 12'h9D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9D8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b110, 12'h9D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b110, 12'h9DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b110, 12'h9E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b110, 12'h9E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9E8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b110, 12'h9E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9EC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b110, 12'h9ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b110, 12'h9F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9F4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b110, 12'h9F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9F8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b110, 12'h9F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'h9FC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b110, 12'h9FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA00} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b110, 12'hA01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA04} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b110, 12'hA05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA08} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b110, 12'hA09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA0C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b110, 12'hA0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA10} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b110, 12'hA11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA14} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b110, 12'hA15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA18} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b110, 12'hA19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA1C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b110, 12'hA1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA20} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b110, 12'hA21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA24} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b110, 12'hA25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA28} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b110, 12'hA29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA2C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b110, 12'hA2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA30} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b110, 12'hA31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA34} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b110, 12'hA35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA38} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b110, 12'hA39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA3C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b110, 12'hA3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA40} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b110, 12'hA41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA44} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b110, 12'hA45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA48} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b110, 12'hA49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA4C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b110, 12'hA4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA50} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b110, 12'hA51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA54} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b110, 12'hA55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA58} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b110, 12'hA59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA5C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b110, 12'hA5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA60} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b110, 12'hA61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA64} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b110, 12'hA65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA68} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b110, 12'hA69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA6C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b110, 12'hA6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA70} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b110, 12'hA71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA74} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b110, 12'hA75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b110, 12'hA79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA7C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b110, 12'hA7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA80} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b110, 12'hA81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA84} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b110, 12'hA85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA88} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b110, 12'hA89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA8C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b110, 12'hA8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA90} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b110, 12'hA91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA94} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b110, 12'hA95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA98} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b110, 12'hA99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hA9C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b110, 12'hA9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAA0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b110, 12'hAA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAA4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b110, 12'hAA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAA8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b110, 12'hAA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAAC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b110, 12'hAAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAB0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b110, 12'hAB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAB4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b110, 12'hAB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAB8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b110, 12'hAB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hABC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b110, 12'hABD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAC0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b110, 12'hAC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAC4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b110, 12'hAC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAC8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b110, 12'hAC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hACC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b110, 12'hACD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAD0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b110, 12'hAD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAD4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b110, 12'hAD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAD8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b110, 12'hAD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hADC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b110, 12'hADD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAE0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b110, 12'hAE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAE4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b110, 12'hAE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAE8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b110, 12'hAE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAEC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b110, 12'hAED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAF0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b110, 12'hAF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAF4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b110, 12'hAF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAF8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b110, 12'hAF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hAFC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b110, 12'hAFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB00} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b110, 12'hB01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB04} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b110, 12'hB05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB08} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b110, 12'hB09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB0C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b110, 12'hB0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB10} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b110, 12'hB11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB14} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b110, 12'hB15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB18} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b110, 12'hB19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB1C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b110, 12'hB1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB20} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b110, 12'hB21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB24} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b110, 12'hB25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB28} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b110, 12'hB29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB2C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b110, 12'hB2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB30} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b110, 12'hB31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB34} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b110, 12'hB35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB38} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b110, 12'hB39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB3C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b110, 12'hB3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB40} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b110, 12'hB41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB44} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b110, 12'hB45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB48} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b110, 12'hB49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB4C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b110, 12'hB4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB50} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b110, 12'hB51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB54} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b110, 12'hB55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB58} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b110, 12'hB59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB5C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b110, 12'hB5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB60} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b110, 12'hB61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB64} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b110, 12'hB65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB68} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b110, 12'hB69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB6C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b110, 12'hB6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB70} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b110, 12'hB71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB74} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b110, 12'hB75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB78} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b110, 12'hB79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB7C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b110, 12'hB7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB80} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b110, 12'hB81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB84} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b110, 12'hB85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB88} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b110, 12'hB89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB8C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b110, 12'hB8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB90} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b110, 12'hB91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB94} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b110, 12'hB95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB98} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b110, 12'hB99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hB9C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b110, 12'hB9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBA0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b110, 12'hBA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBA4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b110, 12'hBA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBA8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b110, 12'hBA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBAC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b110, 12'hBAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBB0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b110, 12'hBB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBB4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b110, 12'hBB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBB8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b110, 12'hBB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBBC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b110, 12'hBBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBC0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b110, 12'hBC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBC4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b110, 12'hBC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBC8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b110, 12'hBC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBCC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b110, 12'hBCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBD0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b110, 12'hBD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBD4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b110, 12'hBD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBD8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b110, 12'hBD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBDC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b110, 12'hBDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBE0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b110, 12'hBE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBE4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b110, 12'hBE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBE8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b110, 12'hBE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBEC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b110, 12'hBED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBF0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b110, 12'hBF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBF4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b110, 12'hBF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBF8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b110, 12'hBF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hBFC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b110, 12'hBFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC04} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b110, 12'hC05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC08} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b110, 12'hC09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC0C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b110, 12'hC0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC10} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b110, 12'hC11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC14} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b110, 12'hC15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC18} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b110, 12'hC19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC1C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b110, 12'hC1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC20} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b110, 12'hC21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC24} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b110, 12'hC25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC28} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b110, 12'hC29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC2C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b110, 12'hC2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC30} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b110, 12'hC31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC34} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b110, 12'hC35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC38} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b110, 12'hC39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC3C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b110, 12'hC3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC40} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC44} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b110, 12'hC45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC48} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b110, 12'hC49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC4C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b110, 12'hC4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC50} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b110, 12'hC51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC54} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b110, 12'hC55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC58} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b110, 12'hC59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC5C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b110, 12'hC5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC60} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b110, 12'hC61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC64} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b110, 12'hC65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC68} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b110, 12'hC69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC6C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b110, 12'hC6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC70} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b110, 12'hC71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC74} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b110, 12'hC75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC78} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b110, 12'hC79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC7C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b110, 12'hC7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC80} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b110, 12'hC81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC84} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b110, 12'hC85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC88} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b110, 12'hC89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC8C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b110, 12'hC8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC90} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b110, 12'hC91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC94} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b110, 12'hC95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC98} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b110, 12'hC99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hC9C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b110, 12'hC9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCA0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b110, 12'hCA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCA4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b110, 12'hCA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCA8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b110, 12'hCA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCAC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b110, 12'hCAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCB0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b110, 12'hCB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCB4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b110, 12'hCB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCB8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b110, 12'hCB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCBC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b110, 12'hCBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCC0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b110, 12'hCC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCC4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b110, 12'hCC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCC8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b110, 12'hCC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCCC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b110, 12'hCCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCD0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b110, 12'hCD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCD4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b110, 12'hCD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCD8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b110, 12'hCD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCDC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b110, 12'hCDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCE0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b110, 12'hCE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCE4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b110, 12'hCE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCE8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b110, 12'hCE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCEC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b110, 12'hCED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCF0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b110, 12'hCF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCF4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b110, 12'hCF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCF8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b110, 12'hCF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hCFC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b110, 12'hCFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD00} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b110, 12'hD01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD04} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b110, 12'hD05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD08} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b110, 12'hD09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD0C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b110, 12'hD0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD10} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b110, 12'hD11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD14} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b110, 12'hD15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD18} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b110, 12'hD19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD1C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b110, 12'hD1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD20} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b110, 12'hD21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD24} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b110, 12'hD25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD28} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b110, 12'hD29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD2C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b110, 12'hD2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD30} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b110, 12'hD31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD34} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b110, 12'hD35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD38} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b110, 12'hD39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD3C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b110, 12'hD3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD40} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b110, 12'hD41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD44} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b110, 12'hD45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD48} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b110, 12'hD49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD4C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b110, 12'hD4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD50} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b110, 12'hD51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD54} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b110, 12'hD55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD58} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b110, 12'hD59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD5C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b110, 12'hD5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD60} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b110, 12'hD61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD64} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b110, 12'hD65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD68} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b110, 12'hD69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD6C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b110, 12'hD6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD70} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b110, 12'hD71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD74} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b110, 12'hD75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD78} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b110, 12'hD79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD7C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b110, 12'hD7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD80} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b110, 12'hD81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD84} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b110, 12'hD85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD88} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b110, 12'hD89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD8C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b110, 12'hD8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD90} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b110, 12'hD91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD94} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b110, 12'hD95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD98} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b110, 12'hD99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hD9C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b110, 12'hD9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDA0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b110, 12'hDA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDA4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b110, 12'hDA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDA8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b110, 12'hDA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDAC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b110, 12'hDAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDB0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b110, 12'hDB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDB4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b110, 12'hDB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDB8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b110, 12'hDB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDBC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b110, 12'hDBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDC0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b110, 12'hDC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDC4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b110, 12'hDC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDC8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b110, 12'hDC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDCC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b110, 12'hDCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDD0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b110, 12'hDD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDD4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b110, 12'hDD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDD8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b110, 12'hDD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDDC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b110, 12'hDDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDE0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b110, 12'hDE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDE4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b110, 12'hDE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDE8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b110, 12'hDE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDEC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b110, 12'hDED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDF0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b110, 12'hDF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDF4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b110, 12'hDF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDF8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b110, 12'hDF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hDFC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b110, 12'hDFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE00} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b110, 12'hE01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE04} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b110, 12'hE05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE08} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b110, 12'hE09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE0C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b110, 12'hE0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE10} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b110, 12'hE11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE14} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b110, 12'hE15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE18} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b110, 12'hE19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE1C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b110, 12'hE1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE20} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b110, 12'hE21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE24} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b110, 12'hE25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE28} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b110, 12'hE29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE2C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b110, 12'hE2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE30} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b110, 12'hE31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE34} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b110, 12'hE35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE38} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b110, 12'hE39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE3C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b110, 12'hE3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE40} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b110, 12'hE41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE44} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b110, 12'hE45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE48} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b110, 12'hE49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE4C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b110, 12'hE4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE50} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b110, 12'hE51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE54} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b110, 12'hE55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE58} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b110, 12'hE59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE5C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b110, 12'hE5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE60} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b110, 12'hE61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE64} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b110, 12'hE65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE68} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b110, 12'hE69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE6C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b110, 12'hE6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE70} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b110, 12'hE71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE74} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b110, 12'hE75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b110, 12'hE79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE7C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b110, 12'hE7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE80} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b110, 12'hE81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE84} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b110, 12'hE85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE88} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b110, 12'hE89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE8C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b110, 12'hE8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE90} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b110, 12'hE91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE94} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b110, 12'hE95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE98} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b110, 12'hE99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hE9C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b110, 12'hE9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEA0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b110, 12'hEA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEA4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b110, 12'hEA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEA8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b110, 12'hEA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEAC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b110, 12'hEAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEB0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b110, 12'hEB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEB4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b110, 12'hEB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEB8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b110, 12'hEB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEBC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b110, 12'hEBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEC0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b110, 12'hEC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEC4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b110, 12'hEC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEC8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b110, 12'hEC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hECC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b110, 12'hECD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hED0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b110, 12'hED1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hED4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b110, 12'hED5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hED8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b110, 12'hED9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEDC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b110, 12'hEDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEE0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b110, 12'hEE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEE4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b110, 12'hEE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEE8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b110, 12'hEE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEEC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b110, 12'hEED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEF0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b110, 12'hEF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEF4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b110, 12'hEF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEF8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b110, 12'hEF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hEFC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b110, 12'hEFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF00} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b110, 12'hF01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF04} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b110, 12'hF05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF08} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b110, 12'hF09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF0C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b110, 12'hF0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF10} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b110, 12'hF11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF14} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b110, 12'hF15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF18} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b110, 12'hF19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF1C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b110, 12'hF1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF20} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b110, 12'hF21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF24} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b110, 12'hF25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF28} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b110, 12'hF29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF2C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b110, 12'hF2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF30} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b110, 12'hF31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF34} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b110, 12'hF35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF38} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b110, 12'hF39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF3C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b110, 12'hF3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF40} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b110, 12'hF41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF44} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b110, 12'hF45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF48} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b110, 12'hF49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF4C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b110, 12'hF4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF50} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b110, 12'hF51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF54} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b110, 12'hF55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF58} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b110, 12'hF59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF5C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b110, 12'hF5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF60} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b110, 12'hF61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF64} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b110, 12'hF65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF68} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b110, 12'hF69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF6C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b110, 12'hF6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF70} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b110, 12'hF71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF74} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b110, 12'hF75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF78} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b110, 12'hF79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF7C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b110, 12'hF7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF80} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b110, 12'hF81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF84} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b110, 12'hF85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF88} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b110, 12'hF89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF8C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b110, 12'hF8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF90} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b110, 12'hF91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF94} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b110, 12'hF95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF98} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b110, 12'hF99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hF9C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b110, 12'hF9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFA0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b110, 12'hFA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFA4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b110, 12'hFA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFA8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b110, 12'hFA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFAC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b110, 12'hFAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFB0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b110, 12'hFB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFB4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b110, 12'hFB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFB8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b110, 12'hFB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFBC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b110, 12'hFBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFC0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b110, 12'hFC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFC4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b110, 12'hFC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFC8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b110, 12'hFC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFCC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b110, 12'hFCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFD0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b110, 12'hFD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFD4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b110, 12'hFD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFD8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b110, 12'hFD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFDC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b110, 12'hFDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFE0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b110, 12'hFE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFE4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b110, 12'hFE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFE8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b110, 12'hFE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFEC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b110, 12'hFED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFF0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b110, 12'hFF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFF4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b110, 12'hFF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFF8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b110, 12'hFF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b110, 12'hFFC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b110, 12'hFFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h001} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h004} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b111, 12'h005} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h008} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b111, 12'h009} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h00C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b111, 12'h00D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h010} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b111, 12'h011} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h014} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b111, 12'h015} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h018} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b111, 12'h019} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h01C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b111, 12'h01D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h020} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b111, 12'h021} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h024} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b111, 12'h025} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h028} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b111, 12'h029} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h02C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b111, 12'h02D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h030} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b111, 12'h031} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h034} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b111, 12'h035} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h038} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b111, 12'h039} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h03C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b111, 12'h03D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h040} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h041} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h044} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b111, 12'h045} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h048} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b111, 12'h049} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h04C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b111, 12'h04D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h050} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b111, 12'h051} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h054} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b111, 12'h055} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h058} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b111, 12'h059} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h05C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b111, 12'h05D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h060} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b111, 12'h061} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h064} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b111, 12'h065} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h068} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b111, 12'h069} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h06C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b111, 12'h06D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h070} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b111, 12'h071} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h074} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b111, 12'h075} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h078} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b111, 12'h079} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h07C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b111, 12'h07D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h080} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b111, 12'h081} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h084} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b111, 12'h085} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h088} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b111, 12'h089} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h08C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b111, 12'h08D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h090} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b111, 12'h091} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h094} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b111, 12'h095} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h098} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b111, 12'h099} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h09C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b111, 12'h09D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0A0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b111, 12'h0A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0A4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b111, 12'h0A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0A8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b111, 12'h0A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0AC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b111, 12'h0AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0B0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b111, 12'h0B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0B4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b111, 12'h0B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0B8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b111, 12'h0B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0BC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b111, 12'h0BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0C0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b111, 12'h0C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0C4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b111, 12'h0C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0C8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b111, 12'h0C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0CC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b111, 12'h0CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0D0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b111, 12'h0D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0D4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b111, 12'h0D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0D8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b111, 12'h0D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0DC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b111, 12'h0DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0E0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b111, 12'h0E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0E4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b111, 12'h0E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0E8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b111, 12'h0E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0EC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b111, 12'h0ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0F0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b111, 12'h0F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0F4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b111, 12'h0F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b111, 12'h0F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h0FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b111, 12'h0FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h100} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b111, 12'h101} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h104} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b111, 12'h105} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h108} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b111, 12'h109} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h10C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b111, 12'h10D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h110} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b111, 12'h111} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h114} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b111, 12'h115} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h118} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b111, 12'h119} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h11C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b111, 12'h11D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h120} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b111, 12'h121} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h124} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b111, 12'h125} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h128} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b111, 12'h129} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h12C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b111, 12'h12D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h130} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b111, 12'h131} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h134} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b111, 12'h135} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h138} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b111, 12'h139} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h13C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b111, 12'h13D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h140} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b111, 12'h141} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h144} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b111, 12'h145} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h148} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b111, 12'h149} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h14C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b111, 12'h14D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h150} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b111, 12'h151} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h154} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b111, 12'h155} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h158} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b111, 12'h159} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h15C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b111, 12'h15D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h160} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b111, 12'h161} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h164} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b111, 12'h165} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h168} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b111, 12'h169} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h16C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b111, 12'h16D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h170} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b111, 12'h171} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h174} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b111, 12'h175} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h178} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b111, 12'h179} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h17C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b111, 12'h17D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h180} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b111, 12'h181} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h184} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b111, 12'h185} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h188} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b111, 12'h189} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h18C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b111, 12'h18D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h190} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b111, 12'h191} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h194} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b111, 12'h195} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h198} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b111, 12'h199} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h19C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b111, 12'h19D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b111, 12'h1A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b111, 12'h1A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b111, 12'h1A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b111, 12'h1AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b111, 12'h1B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b111, 12'h1B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b111, 12'h1B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b111, 12'h1BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1C0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b111, 12'h1C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b111, 12'h1C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1C8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b111, 12'h1C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1CC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b111, 12'h1CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1D0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b111, 12'h1D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1D4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b111, 12'h1D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1D8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b111, 12'h1D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b111, 12'h1DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b111, 12'h1E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b111, 12'h1E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1E8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b111, 12'h1E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1EC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b111, 12'h1ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b111, 12'h1F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1F4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b111, 12'h1F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1F8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b111, 12'h1F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h1FC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b111, 12'h1FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h200} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b111, 12'h201} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h204} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b111, 12'h205} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h208} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b111, 12'h209} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h20C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b111, 12'h20D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h210} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b111, 12'h211} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h214} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b111, 12'h215} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h218} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b111, 12'h219} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h21C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b111, 12'h21D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h220} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b111, 12'h221} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h224} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b111, 12'h225} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h228} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b111, 12'h229} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h22C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b111, 12'h22D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h230} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b111, 12'h231} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h234} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b111, 12'h235} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h238} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b111, 12'h239} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h23C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b111, 12'h23D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h240} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b111, 12'h241} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h244} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b111, 12'h245} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h248} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b111, 12'h249} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h24C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b111, 12'h24D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h250} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b111, 12'h251} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h254} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b111, 12'h255} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h258} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b111, 12'h259} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h25C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b111, 12'h25D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h260} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b111, 12'h261} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h264} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b111, 12'h265} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h268} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b111, 12'h269} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h26C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b111, 12'h26D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h270} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b111, 12'h271} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h274} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b111, 12'h275} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h278} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b111, 12'h279} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h27C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b111, 12'h27D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h280} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b111, 12'h281} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h284} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b111, 12'h285} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h288} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b111, 12'h289} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h28C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b111, 12'h28D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h290} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b111, 12'h291} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h294} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b111, 12'h295} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h298} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b111, 12'h299} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h29C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b111, 12'h29D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2A0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b111, 12'h2A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2A4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b111, 12'h2A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2A8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b111, 12'h2A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2AC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b111, 12'h2AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2B0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b111, 12'h2B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2B4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b111, 12'h2B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2B8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b111, 12'h2B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2BC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b111, 12'h2BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2C0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b111, 12'h2C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2C4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b111, 12'h2C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2C8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b111, 12'h2C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2CC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b111, 12'h2CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2D0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b111, 12'h2D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2D4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b111, 12'h2D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2D8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b111, 12'h2D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2DC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b111, 12'h2DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2E0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b111, 12'h2E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2E4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b111, 12'h2E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2E8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b111, 12'h2E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2EC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b111, 12'h2ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2F0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b111, 12'h2F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2F4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b111, 12'h2F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2F8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b111, 12'h2F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h2FC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b111, 12'h2FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h300} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b111, 12'h301} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h304} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b111, 12'h305} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h308} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b111, 12'h309} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h30C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b111, 12'h30D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h310} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b111, 12'h311} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h314} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b111, 12'h315} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h318} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b111, 12'h319} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h31C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b111, 12'h31D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h320} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b111, 12'h321} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h324} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b111, 12'h325} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h328} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b111, 12'h329} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h32C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b111, 12'h32D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h330} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b111, 12'h331} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h334} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b111, 12'h335} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h338} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b111, 12'h339} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h33C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b111, 12'h33D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h340} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b111, 12'h341} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h344} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b111, 12'h345} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h348} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b111, 12'h349} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h34C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b111, 12'h34D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h350} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b111, 12'h351} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h354} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b111, 12'h355} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h358} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b111, 12'h359} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h35C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b111, 12'h35D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h360} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b111, 12'h361} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h364} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b111, 12'h365} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h368} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b111, 12'h369} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h36C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b111, 12'h36D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h370} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b111, 12'h371} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h374} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b111, 12'h375} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h378} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b111, 12'h379} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h37C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b111, 12'h37D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h380} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b111, 12'h381} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h384} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b111, 12'h385} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h388} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b111, 12'h389} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h38C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b111, 12'h38D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h390} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b111, 12'h391} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h394} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b111, 12'h395} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h398} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b111, 12'h399} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h39C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b111, 12'h39D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3A0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b111, 12'h3A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3A4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b111, 12'h3A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3A8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b111, 12'h3A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3AC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b111, 12'h3AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3B0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b111, 12'h3B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3B4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b111, 12'h3B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3B8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b111, 12'h3B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3BC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b111, 12'h3BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3C0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b111, 12'h3C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3C4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b111, 12'h3C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3C8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b111, 12'h3C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3CC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b111, 12'h3CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3D0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b111, 12'h3D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3D4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b111, 12'h3D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3D8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b111, 12'h3D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3DC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b111, 12'h3DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3E0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b111, 12'h3E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3E4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b111, 12'h3E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3E8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b111, 12'h3E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3EC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b111, 12'h3ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3F0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b111, 12'h3F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3F4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b111, 12'h3F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3F8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b111, 12'h3F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h3FC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b111, 12'h3FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h401} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h404} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b111, 12'h405} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h408} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b111, 12'h409} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h40C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b111, 12'h40D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h410} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b111, 12'h411} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h414} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b111, 12'h415} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h418} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b111, 12'h419} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h41C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b111, 12'h41D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h420} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b111, 12'h421} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h424} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b111, 12'h425} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h428} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b111, 12'h429} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h42C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b111, 12'h42D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h430} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b111, 12'h431} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h434} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b111, 12'h435} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h438} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b111, 12'h439} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h43C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b111, 12'h43D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h440} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h441} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h444} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b111, 12'h445} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h448} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b111, 12'h449} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h44C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b111, 12'h44D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h450} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b111, 12'h451} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h454} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b111, 12'h455} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h458} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b111, 12'h459} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h45C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b111, 12'h45D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h460} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b111, 12'h461} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h464} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b111, 12'h465} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h468} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b111, 12'h469} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h46C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b111, 12'h46D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h470} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b111, 12'h471} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h474} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b111, 12'h475} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h478} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b111, 12'h479} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h47C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b111, 12'h47D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h480} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b111, 12'h481} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h484} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b111, 12'h485} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h488} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b111, 12'h489} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h48C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b111, 12'h48D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h490} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b111, 12'h491} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h494} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b111, 12'h495} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h498} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b111, 12'h499} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h49C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b111, 12'h49D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4A0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b111, 12'h4A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4A4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b111, 12'h4A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4A8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b111, 12'h4A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4AC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b111, 12'h4AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4B0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b111, 12'h4B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4B4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b111, 12'h4B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4B8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b111, 12'h4B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4BC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b111, 12'h4BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4C0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b111, 12'h4C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4C4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b111, 12'h4C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4C8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b111, 12'h4C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4CC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b111, 12'h4CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4D0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b111, 12'h4D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4D4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b111, 12'h4D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4D8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b111, 12'h4D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4DC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b111, 12'h4DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4E0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b111, 12'h4E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4E4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b111, 12'h4E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4E8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b111, 12'h4E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4EC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b111, 12'h4ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4F0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b111, 12'h4F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4F4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b111, 12'h4F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b111, 12'h4F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h4FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b111, 12'h4FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h500} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b111, 12'h501} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h504} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b111, 12'h505} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h508} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b111, 12'h509} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h50C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b111, 12'h50D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h510} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b111, 12'h511} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h514} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b111, 12'h515} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h518} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b111, 12'h519} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h51C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b111, 12'h51D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h520} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b111, 12'h521} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h524} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b111, 12'h525} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h528} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b111, 12'h529} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h52C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b111, 12'h52D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h530} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b111, 12'h531} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h534} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b111, 12'h535} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h538} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b111, 12'h539} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h53C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b111, 12'h53D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h540} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b111, 12'h541} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h544} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b111, 12'h545} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h548} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b111, 12'h549} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h54C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b111, 12'h54D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h550} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b111, 12'h551} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h554} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b111, 12'h555} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h558} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b111, 12'h559} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h55C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b111, 12'h55D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h560} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b111, 12'h561} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h564} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b111, 12'h565} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h568} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b111, 12'h569} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h56C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b111, 12'h56D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h570} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b111, 12'h571} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h574} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b111, 12'h575} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h578} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b111, 12'h579} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h57C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b111, 12'h57D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h580} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b111, 12'h581} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h584} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b111, 12'h585} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h588} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b111, 12'h589} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h58C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b111, 12'h58D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h590} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b111, 12'h591} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h594} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b111, 12'h595} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h598} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b111, 12'h599} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h59C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b111, 12'h59D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b111, 12'h5A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b111, 12'h5A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b111, 12'h5A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b111, 12'h5AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b111, 12'h5B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b111, 12'h5B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b111, 12'h5B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b111, 12'h5BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5C0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b111, 12'h5C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b111, 12'h5C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5C8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b111, 12'h5C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5CC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b111, 12'h5CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5D0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b111, 12'h5D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5D4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b111, 12'h5D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5D8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b111, 12'h5D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b111, 12'h5DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b111, 12'h5E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b111, 12'h5E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5E8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b111, 12'h5E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5EC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b111, 12'h5ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b111, 12'h5F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5F4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b111, 12'h5F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5F8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b111, 12'h5F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h5FC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b111, 12'h5FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h600} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b111, 12'h601} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h604} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b111, 12'h605} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h608} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b111, 12'h609} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h60C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b111, 12'h60D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h610} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b111, 12'h611} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h614} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b111, 12'h615} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h618} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b111, 12'h619} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h61C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b111, 12'h61D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h620} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b111, 12'h621} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h624} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b111, 12'h625} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h628} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b111, 12'h629} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h62C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b111, 12'h62D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h630} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b111, 12'h631} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h634} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b111, 12'h635} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h638} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b111, 12'h639} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h63C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b111, 12'h63D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h640} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b111, 12'h641} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h644} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b111, 12'h645} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h648} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b111, 12'h649} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h64C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b111, 12'h64D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h650} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b111, 12'h651} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h654} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b111, 12'h655} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h658} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b111, 12'h659} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h65C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b111, 12'h65D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h660} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b111, 12'h661} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h664} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b111, 12'h665} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h668} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b111, 12'h669} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h66C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b111, 12'h66D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h670} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b111, 12'h671} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h674} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b111, 12'h675} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h678} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b111, 12'h679} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h67C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b111, 12'h67D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h680} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b111, 12'h681} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h684} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b111, 12'h685} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h688} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b111, 12'h689} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h68C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b111, 12'h68D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h690} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b111, 12'h691} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h694} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b111, 12'h695} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h698} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b111, 12'h699} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h69C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b111, 12'h69D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6A0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b111, 12'h6A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6A4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b111, 12'h6A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6A8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b111, 12'h6A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6AC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b111, 12'h6AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6B0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b111, 12'h6B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6B4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b111, 12'h6B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6B8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b111, 12'h6B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6BC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b111, 12'h6BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6C0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b111, 12'h6C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6C4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b111, 12'h6C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6C8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b111, 12'h6C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6CC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b111, 12'h6CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6D0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b111, 12'h6D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6D4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b111, 12'h6D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6D8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b111, 12'h6D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6DC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b111, 12'h6DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6E0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b111, 12'h6E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6E4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b111, 12'h6E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6E8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b111, 12'h6E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6EC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b111, 12'h6ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6F0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b111, 12'h6F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6F4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b111, 12'h6F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6F8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b111, 12'h6F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h6FC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b111, 12'h6FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h700} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b111, 12'h701} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h704} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b111, 12'h705} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h708} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b111, 12'h709} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h70C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b111, 12'h70D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h710} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b111, 12'h711} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h714} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b111, 12'h715} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h718} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b111, 12'h719} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h71C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b111, 12'h71D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h720} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b111, 12'h721} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h724} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b111, 12'h725} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h728} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b111, 12'h729} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h72C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b111, 12'h72D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h730} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b111, 12'h731} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h734} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b111, 12'h735} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h738} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b111, 12'h739} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h73C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b111, 12'h73D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h740} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b111, 12'h741} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h744} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b111, 12'h745} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h748} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b111, 12'h749} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h74C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b111, 12'h74D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h750} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b111, 12'h751} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h754} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b111, 12'h755} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h758} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b111, 12'h759} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h75C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b111, 12'h75D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h760} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b111, 12'h761} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h764} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b111, 12'h765} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h768} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b111, 12'h769} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h76C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b111, 12'h76D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h770} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b111, 12'h771} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h774} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b111, 12'h775} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h778} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b111, 12'h779} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h77C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b111, 12'h77D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h780} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b111, 12'h781} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h784} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b111, 12'h785} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h788} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b111, 12'h789} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h78C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b111, 12'h78D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h790} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b111, 12'h791} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h794} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b111, 12'h795} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h798} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b111, 12'h799} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h79C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b111, 12'h79D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7A0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b111, 12'h7A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7A4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b111, 12'h7A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7A8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b111, 12'h7A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7AC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b111, 12'h7AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7B0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b111, 12'h7B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7B4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b111, 12'h7B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7B8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b111, 12'h7B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7BC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b111, 12'h7BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7C0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b111, 12'h7C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7C4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b111, 12'h7C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7C8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b111, 12'h7C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7CC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b111, 12'h7CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7D0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b111, 12'h7D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7D4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b111, 12'h7D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7D8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b111, 12'h7D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7DC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b111, 12'h7DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7E0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b111, 12'h7E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7E4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b111, 12'h7E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7E8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b111, 12'h7E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7EC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b111, 12'h7ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7F0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b111, 12'h7F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7F4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b111, 12'h7F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7F8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b111, 12'h7F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h7FC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b111, 12'h7FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h801} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h804} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b111, 12'h805} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h808} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b111, 12'h809} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h80C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b111, 12'h80D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h810} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b111, 12'h811} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h814} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b111, 12'h815} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h818} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b111, 12'h819} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h81C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b111, 12'h81D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h820} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b111, 12'h821} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h824} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b111, 12'h825} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h828} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b111, 12'h829} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h82C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b111, 12'h82D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h830} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b111, 12'h831} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h834} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b111, 12'h835} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h838} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b111, 12'h839} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h83C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b111, 12'h83D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h840} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h841} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h844} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b111, 12'h845} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h848} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b111, 12'h849} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h84C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b111, 12'h84D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h850} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b111, 12'h851} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h854} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b111, 12'h855} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h858} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b111, 12'h859} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h85C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b111, 12'h85D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h860} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b111, 12'h861} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h864} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b111, 12'h865} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h868} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b111, 12'h869} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h86C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b111, 12'h86D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h870} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b111, 12'h871} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h874} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b111, 12'h875} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h878} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b111, 12'h879} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h87C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b111, 12'h87D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h880} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b111, 12'h881} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h884} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b111, 12'h885} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h888} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b111, 12'h889} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h88C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b111, 12'h88D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h890} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b111, 12'h891} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h894} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b111, 12'h895} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h898} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b111, 12'h899} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h89C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b111, 12'h89D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8A0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b111, 12'h8A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8A4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b111, 12'h8A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8A8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b111, 12'h8A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8AC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b111, 12'h8AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8B0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b111, 12'h8B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8B4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b111, 12'h8B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8B8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b111, 12'h8B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8BC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b111, 12'h8BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8C0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b111, 12'h8C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8C4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b111, 12'h8C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8C8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b111, 12'h8C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8CC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b111, 12'h8CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8D0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b111, 12'h8D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8D4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b111, 12'h8D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8D8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b111, 12'h8D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8DC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b111, 12'h8DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8E0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b111, 12'h8E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8E4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b111, 12'h8E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8E8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b111, 12'h8E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8EC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b111, 12'h8ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8F0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b111, 12'h8F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8F4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b111, 12'h8F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8F8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b111, 12'h8F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h8FC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b111, 12'h8FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h900} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b111, 12'h901} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h904} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b111, 12'h905} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h908} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b111, 12'h909} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h90C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b111, 12'h90D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h910} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b111, 12'h911} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h914} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b111, 12'h915} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h918} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b111, 12'h919} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h91C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b111, 12'h91D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h920} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b111, 12'h921} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h924} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b111, 12'h925} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h928} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b111, 12'h929} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h92C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b111, 12'h92D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h930} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b111, 12'h931} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h934} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b111, 12'h935} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h938} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b111, 12'h939} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h93C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b111, 12'h93D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h940} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b111, 12'h941} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h944} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b111, 12'h945} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h948} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b111, 12'h949} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h94C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b111, 12'h94D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h950} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b111, 12'h951} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h954} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b111, 12'h955} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h958} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b111, 12'h959} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h95C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b111, 12'h95D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h960} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b111, 12'h961} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h964} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b111, 12'h965} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h968} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b111, 12'h969} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h96C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b111, 12'h96D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h970} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b111, 12'h971} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h974} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b111, 12'h975} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h978} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b111, 12'h979} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h97C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b111, 12'h97D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h980} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b111, 12'h981} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h984} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b111, 12'h985} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h988} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b111, 12'h989} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h98C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b111, 12'h98D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h990} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b111, 12'h991} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h994} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b111, 12'h995} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h998} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b111, 12'h999} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h99C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b111, 12'h99D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9A0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b111, 12'h9A1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9A4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b111, 12'h9A5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9A8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b111, 12'h9A9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9AC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b111, 12'h9AD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9B0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b111, 12'h9B1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9B4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b111, 12'h9B5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9B8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b111, 12'h9B9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9BC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b111, 12'h9BD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9C0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b111, 12'h9C1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9C4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b111, 12'h9C5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9C8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b111, 12'h9C9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9CC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b111, 12'h9CD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9D0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b111, 12'h9D1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9D4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b111, 12'h9D5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9D8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b111, 12'h9D9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9DC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b111, 12'h9DD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9E0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b111, 12'h9E1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9E4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b111, 12'h9E5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9E8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b111, 12'h9E9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9EC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b111, 12'h9ED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9F0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b111, 12'h9F1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9F4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b111, 12'h9F5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9F8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b111, 12'h9F9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'h9FC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b111, 12'h9FD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA00} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b111, 12'hA01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA04} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b111, 12'hA05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA08} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b111, 12'hA09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA0C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b111, 12'hA0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA10} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b111, 12'hA11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA14} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b111, 12'hA15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA18} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b111, 12'hA19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA1C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b111, 12'hA1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA20} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b111, 12'hA21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA24} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b111, 12'hA25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA28} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b111, 12'hA29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA2C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b111, 12'hA2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA30} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b111, 12'hA31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA34} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b111, 12'hA35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA38} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b111, 12'hA39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA3C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b111, 12'hA3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA40} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b111, 12'hA41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA44} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b111, 12'hA45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA48} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b111, 12'hA49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA4C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b111, 12'hA4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA50} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b111, 12'hA51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA54} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b111, 12'hA55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA58} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b111, 12'hA59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA5C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b111, 12'hA5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA60} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b111, 12'hA61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA64} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b111, 12'hA65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA68} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b111, 12'hA69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA6C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b111, 12'hA6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA70} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b111, 12'hA71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA74} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b111, 12'hA75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b111, 12'hA79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA7C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b111, 12'hA7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA80} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b111, 12'hA81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA84} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b111, 12'hA85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA88} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b111, 12'hA89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA8C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b111, 12'hA8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA90} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b111, 12'hA91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA94} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b111, 12'hA95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA98} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b111, 12'hA99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hA9C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b111, 12'hA9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAA0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b111, 12'hAA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAA4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b111, 12'hAA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAA8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b111, 12'hAA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAAC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b111, 12'hAAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAB0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b111, 12'hAB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAB4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b111, 12'hAB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAB8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b111, 12'hAB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hABC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b111, 12'hABD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAC0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b111, 12'hAC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAC4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b111, 12'hAC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAC8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b111, 12'hAC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hACC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b111, 12'hACD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAD0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b111, 12'hAD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAD4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b111, 12'hAD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAD8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b111, 12'hAD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hADC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b111, 12'hADD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAE0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b111, 12'hAE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAE4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b111, 12'hAE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAE8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b111, 12'hAE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAEC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b111, 12'hAED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAF0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b111, 12'hAF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAF4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b111, 12'hAF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAF8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b111, 12'hAF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hAFC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b111, 12'hAFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB00} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b111, 12'hB01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB04} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b111, 12'hB05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB08} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b111, 12'hB09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB0C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b111, 12'hB0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB10} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b111, 12'hB11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB14} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b111, 12'hB15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB18} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b111, 12'hB19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB1C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b111, 12'hB1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB20} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b111, 12'hB21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB24} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b111, 12'hB25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB28} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b111, 12'hB29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB2C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b111, 12'hB2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB30} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b111, 12'hB31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB34} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b111, 12'hB35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB38} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b111, 12'hB39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB3C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b111, 12'hB3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB40} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b111, 12'hB41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB44} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b111, 12'hB45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB48} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b111, 12'hB49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB4C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b111, 12'hB4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB50} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b111, 12'hB51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB54} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b111, 12'hB55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB58} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b111, 12'hB59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB5C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b111, 12'hB5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB60} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b111, 12'hB61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB64} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b111, 12'hB65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB68} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b111, 12'hB69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB6C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b111, 12'hB6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB70} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b111, 12'hB71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB74} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b111, 12'hB75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB78} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b111, 12'hB79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB7C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b111, 12'hB7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB80} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b111, 12'hB81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB84} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b111, 12'hB85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB88} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b111, 12'hB89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB8C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b111, 12'hB8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB90} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b111, 12'hB91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB94} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b111, 12'hB95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB98} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b111, 12'hB99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hB9C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b111, 12'hB9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBA0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b111, 12'hBA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBA4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b111, 12'hBA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBA8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b111, 12'hBA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBAC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b111, 12'hBAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBB0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b111, 12'hBB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBB4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b111, 12'hBB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBB8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b111, 12'hBB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBBC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b111, 12'hBBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBC0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b111, 12'hBC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBC4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b111, 12'hBC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBC8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b111, 12'hBC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBCC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b111, 12'hBCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBD0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b111, 12'hBD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBD4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b111, 12'hBD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBD8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b111, 12'hBD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBDC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b111, 12'hBDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBE0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b111, 12'hBE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBE4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b111, 12'hBE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBE8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b111, 12'hBE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBEC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b111, 12'hBED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBF0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b111, 12'hBF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBF4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b111, 12'hBF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBF8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b111, 12'hBF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hBFC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b111, 12'hBFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC04} : s_CHIP_23B_45132_reg = 8'h01;
         {3'b111, 12'hC05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC08} : s_CHIP_23B_45132_reg = 8'h02;
         {3'b111, 12'hC09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC0C} : s_CHIP_23B_45132_reg = 8'h03;
         {3'b111, 12'hC0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC10} : s_CHIP_23B_45132_reg = 8'h04;
         {3'b111, 12'hC11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC14} : s_CHIP_23B_45132_reg = 8'h05;
         {3'b111, 12'hC15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC18} : s_CHIP_23B_45132_reg = 8'h06;
         {3'b111, 12'hC19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC1C} : s_CHIP_23B_45132_reg = 8'h07;
         {3'b111, 12'hC1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC20} : s_CHIP_23B_45132_reg = 8'h08;
         {3'b111, 12'hC21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC24} : s_CHIP_23B_45132_reg = 8'h09;
         {3'b111, 12'hC25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC28} : s_CHIP_23B_45132_reg = 8'h0A;
         {3'b111, 12'hC29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC2C} : s_CHIP_23B_45132_reg = 8'h0B;
         {3'b111, 12'hC2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC30} : s_CHIP_23B_45132_reg = 8'h0C;
         {3'b111, 12'hC31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC34} : s_CHIP_23B_45132_reg = 8'h0D;
         {3'b111, 12'hC35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC38} : s_CHIP_23B_45132_reg = 8'h0E;
         {3'b111, 12'hC39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC3C} : s_CHIP_23B_45132_reg = 8'h0F;
         {3'b111, 12'hC3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC40} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC44} : s_CHIP_23B_45132_reg = 8'h11;
         {3'b111, 12'hC45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC48} : s_CHIP_23B_45132_reg = 8'h12;
         {3'b111, 12'hC49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC4C} : s_CHIP_23B_45132_reg = 8'h13;
         {3'b111, 12'hC4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC50} : s_CHIP_23B_45132_reg = 8'h14;
         {3'b111, 12'hC51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC54} : s_CHIP_23B_45132_reg = 8'h15;
         {3'b111, 12'hC55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC58} : s_CHIP_23B_45132_reg = 8'h16;
         {3'b111, 12'hC59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC5C} : s_CHIP_23B_45132_reg = 8'h17;
         {3'b111, 12'hC5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC60} : s_CHIP_23B_45132_reg = 8'h18;
         {3'b111, 12'hC61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC64} : s_CHIP_23B_45132_reg = 8'h19;
         {3'b111, 12'hC65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC68} : s_CHIP_23B_45132_reg = 8'h1A;
         {3'b111, 12'hC69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC6C} : s_CHIP_23B_45132_reg = 8'h1B;
         {3'b111, 12'hC6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC70} : s_CHIP_23B_45132_reg = 8'h1C;
         {3'b111, 12'hC71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC74} : s_CHIP_23B_45132_reg = 8'h1D;
         {3'b111, 12'hC75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC78} : s_CHIP_23B_45132_reg = 8'h1E;
         {3'b111, 12'hC79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC7C} : s_CHIP_23B_45132_reg = 8'h1F;
         {3'b111, 12'hC7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC80} : s_CHIP_23B_45132_reg = 8'h20;
         {3'b111, 12'hC81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC84} : s_CHIP_23B_45132_reg = 8'h21;
         {3'b111, 12'hC85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC88} : s_CHIP_23B_45132_reg = 8'h22;
         {3'b111, 12'hC89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC8C} : s_CHIP_23B_45132_reg = 8'h23;
         {3'b111, 12'hC8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC90} : s_CHIP_23B_45132_reg = 8'h24;
         {3'b111, 12'hC91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC94} : s_CHIP_23B_45132_reg = 8'h25;
         {3'b111, 12'hC95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC98} : s_CHIP_23B_45132_reg = 8'h26;
         {3'b111, 12'hC99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hC9C} : s_CHIP_23B_45132_reg = 8'h27;
         {3'b111, 12'hC9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCA0} : s_CHIP_23B_45132_reg = 8'h28;
         {3'b111, 12'hCA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCA4} : s_CHIP_23B_45132_reg = 8'h29;
         {3'b111, 12'hCA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCA8} : s_CHIP_23B_45132_reg = 8'h2A;
         {3'b111, 12'hCA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCAC} : s_CHIP_23B_45132_reg = 8'h2B;
         {3'b111, 12'hCAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCB0} : s_CHIP_23B_45132_reg = 8'h2C;
         {3'b111, 12'hCB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCB4} : s_CHIP_23B_45132_reg = 8'h2D;
         {3'b111, 12'hCB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCB8} : s_CHIP_23B_45132_reg = 8'h2E;
         {3'b111, 12'hCB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCBC} : s_CHIP_23B_45132_reg = 8'h2F;
         {3'b111, 12'hCBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCC0} : s_CHIP_23B_45132_reg = 8'h30;
         {3'b111, 12'hCC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCC4} : s_CHIP_23B_45132_reg = 8'h31;
         {3'b111, 12'hCC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCC8} : s_CHIP_23B_45132_reg = 8'h32;
         {3'b111, 12'hCC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCCC} : s_CHIP_23B_45132_reg = 8'h33;
         {3'b111, 12'hCCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCD0} : s_CHIP_23B_45132_reg = 8'h34;
         {3'b111, 12'hCD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCD4} : s_CHIP_23B_45132_reg = 8'h35;
         {3'b111, 12'hCD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCD8} : s_CHIP_23B_45132_reg = 8'h36;
         {3'b111, 12'hCD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCDC} : s_CHIP_23B_45132_reg = 8'h37;
         {3'b111, 12'hCDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCE0} : s_CHIP_23B_45132_reg = 8'h38;
         {3'b111, 12'hCE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCE4} : s_CHIP_23B_45132_reg = 8'h39;
         {3'b111, 12'hCE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCE8} : s_CHIP_23B_45132_reg = 8'h3A;
         {3'b111, 12'hCE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCEC} : s_CHIP_23B_45132_reg = 8'h3B;
         {3'b111, 12'hCED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCF0} : s_CHIP_23B_45132_reg = 8'h3C;
         {3'b111, 12'hCF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCF4} : s_CHIP_23B_45132_reg = 8'h3D;
         {3'b111, 12'hCF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCF8} : s_CHIP_23B_45132_reg = 8'h3E;
         {3'b111, 12'hCF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hCFC} : s_CHIP_23B_45132_reg = 8'h3F;
         {3'b111, 12'hCFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD00} : s_CHIP_23B_45132_reg = 8'h40;
         {3'b111, 12'hD01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD04} : s_CHIP_23B_45132_reg = 8'h41;
         {3'b111, 12'hD05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD08} : s_CHIP_23B_45132_reg = 8'h42;
         {3'b111, 12'hD09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD0C} : s_CHIP_23B_45132_reg = 8'h43;
         {3'b111, 12'hD0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD10} : s_CHIP_23B_45132_reg = 8'h44;
         {3'b111, 12'hD11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD14} : s_CHIP_23B_45132_reg = 8'h45;
         {3'b111, 12'hD15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD18} : s_CHIP_23B_45132_reg = 8'h46;
         {3'b111, 12'hD19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD1C} : s_CHIP_23B_45132_reg = 8'h47;
         {3'b111, 12'hD1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD20} : s_CHIP_23B_45132_reg = 8'h48;
         {3'b111, 12'hD21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD24} : s_CHIP_23B_45132_reg = 8'h49;
         {3'b111, 12'hD25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD28} : s_CHIP_23B_45132_reg = 8'h4A;
         {3'b111, 12'hD29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD2C} : s_CHIP_23B_45132_reg = 8'h4B;
         {3'b111, 12'hD2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD30} : s_CHIP_23B_45132_reg = 8'h4C;
         {3'b111, 12'hD31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD34} : s_CHIP_23B_45132_reg = 8'h4D;
         {3'b111, 12'hD35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD38} : s_CHIP_23B_45132_reg = 8'h4E;
         {3'b111, 12'hD39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD3C} : s_CHIP_23B_45132_reg = 8'h4F;
         {3'b111, 12'hD3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD40} : s_CHIP_23B_45132_reg = 8'h50;
         {3'b111, 12'hD41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD44} : s_CHIP_23B_45132_reg = 8'h51;
         {3'b111, 12'hD45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD48} : s_CHIP_23B_45132_reg = 8'h52;
         {3'b111, 12'hD49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD4C} : s_CHIP_23B_45132_reg = 8'h53;
         {3'b111, 12'hD4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD50} : s_CHIP_23B_45132_reg = 8'h54;
         {3'b111, 12'hD51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD54} : s_CHIP_23B_45132_reg = 8'h55;
         {3'b111, 12'hD55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD58} : s_CHIP_23B_45132_reg = 8'h56;
         {3'b111, 12'hD59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD5C} : s_CHIP_23B_45132_reg = 8'h57;
         {3'b111, 12'hD5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD60} : s_CHIP_23B_45132_reg = 8'h58;
         {3'b111, 12'hD61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD64} : s_CHIP_23B_45132_reg = 8'h59;
         {3'b111, 12'hD65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD68} : s_CHIP_23B_45132_reg = 8'h5A;
         {3'b111, 12'hD69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD6C} : s_CHIP_23B_45132_reg = 8'h5B;
         {3'b111, 12'hD6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD70} : s_CHIP_23B_45132_reg = 8'h5C;
         {3'b111, 12'hD71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD74} : s_CHIP_23B_45132_reg = 8'h5D;
         {3'b111, 12'hD75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD78} : s_CHIP_23B_45132_reg = 8'h5E;
         {3'b111, 12'hD79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD7C} : s_CHIP_23B_45132_reg = 8'h5F;
         {3'b111, 12'hD7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD80} : s_CHIP_23B_45132_reg = 8'h60;
         {3'b111, 12'hD81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD84} : s_CHIP_23B_45132_reg = 8'h61;
         {3'b111, 12'hD85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD88} : s_CHIP_23B_45132_reg = 8'h62;
         {3'b111, 12'hD89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD8C} : s_CHIP_23B_45132_reg = 8'h63;
         {3'b111, 12'hD8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD90} : s_CHIP_23B_45132_reg = 8'h64;
         {3'b111, 12'hD91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD94} : s_CHIP_23B_45132_reg = 8'h65;
         {3'b111, 12'hD95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD98} : s_CHIP_23B_45132_reg = 8'h66;
         {3'b111, 12'hD99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hD9C} : s_CHIP_23B_45132_reg = 8'h67;
         {3'b111, 12'hD9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDA0} : s_CHIP_23B_45132_reg = 8'h68;
         {3'b111, 12'hDA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDA4} : s_CHIP_23B_45132_reg = 8'h69;
         {3'b111, 12'hDA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDA8} : s_CHIP_23B_45132_reg = 8'h6A;
         {3'b111, 12'hDA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDAC} : s_CHIP_23B_45132_reg = 8'h6B;
         {3'b111, 12'hDAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDB0} : s_CHIP_23B_45132_reg = 8'h6C;
         {3'b111, 12'hDB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDB4} : s_CHIP_23B_45132_reg = 8'h6D;
         {3'b111, 12'hDB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDB8} : s_CHIP_23B_45132_reg = 8'h6E;
         {3'b111, 12'hDB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDBC} : s_CHIP_23B_45132_reg = 8'h6F;
         {3'b111, 12'hDBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDC0} : s_CHIP_23B_45132_reg = 8'h70;
         {3'b111, 12'hDC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDC4} : s_CHIP_23B_45132_reg = 8'h71;
         {3'b111, 12'hDC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDC8} : s_CHIP_23B_45132_reg = 8'h72;
         {3'b111, 12'hDC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDCC} : s_CHIP_23B_45132_reg = 8'h73;
         {3'b111, 12'hDCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDD0} : s_CHIP_23B_45132_reg = 8'h74;
         {3'b111, 12'hDD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDD4} : s_CHIP_23B_45132_reg = 8'h75;
         {3'b111, 12'hDD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDD8} : s_CHIP_23B_45132_reg = 8'h76;
         {3'b111, 12'hDD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDDC} : s_CHIP_23B_45132_reg = 8'h77;
         {3'b111, 12'hDDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDE0} : s_CHIP_23B_45132_reg = 8'h78;
         {3'b111, 12'hDE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDE4} : s_CHIP_23B_45132_reg = 8'h79;
         {3'b111, 12'hDE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDE8} : s_CHIP_23B_45132_reg = 8'h7A;
         {3'b111, 12'hDE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDEC} : s_CHIP_23B_45132_reg = 8'h7B;
         {3'b111, 12'hDED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDF0} : s_CHIP_23B_45132_reg = 8'h7C;
         {3'b111, 12'hDF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDF4} : s_CHIP_23B_45132_reg = 8'h7D;
         {3'b111, 12'hDF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDF8} : s_CHIP_23B_45132_reg = 8'h7E;
         {3'b111, 12'hDF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hDFC} : s_CHIP_23B_45132_reg = 8'h7F;
         {3'b111, 12'hDFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE00} : s_CHIP_23B_45132_reg = 8'h80;
         {3'b111, 12'hE01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE04} : s_CHIP_23B_45132_reg = 8'h81;
         {3'b111, 12'hE05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE08} : s_CHIP_23B_45132_reg = 8'h82;
         {3'b111, 12'hE09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE0C} : s_CHIP_23B_45132_reg = 8'h83;
         {3'b111, 12'hE0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE10} : s_CHIP_23B_45132_reg = 8'h84;
         {3'b111, 12'hE11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE14} : s_CHIP_23B_45132_reg = 8'h85;
         {3'b111, 12'hE15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE18} : s_CHIP_23B_45132_reg = 8'h86;
         {3'b111, 12'hE19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE1C} : s_CHIP_23B_45132_reg = 8'h87;
         {3'b111, 12'hE1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE20} : s_CHIP_23B_45132_reg = 8'h88;
         {3'b111, 12'hE21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE24} : s_CHIP_23B_45132_reg = 8'h89;
         {3'b111, 12'hE25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE28} : s_CHIP_23B_45132_reg = 8'h8A;
         {3'b111, 12'hE29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE2C} : s_CHIP_23B_45132_reg = 8'h8B;
         {3'b111, 12'hE2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE30} : s_CHIP_23B_45132_reg = 8'h8C;
         {3'b111, 12'hE31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE34} : s_CHIP_23B_45132_reg = 8'h8D;
         {3'b111, 12'hE35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE38} : s_CHIP_23B_45132_reg = 8'h8E;
         {3'b111, 12'hE39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE3C} : s_CHIP_23B_45132_reg = 8'h8F;
         {3'b111, 12'hE3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE40} : s_CHIP_23B_45132_reg = 8'h90;
         {3'b111, 12'hE41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE44} : s_CHIP_23B_45132_reg = 8'h91;
         {3'b111, 12'hE45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE48} : s_CHIP_23B_45132_reg = 8'h92;
         {3'b111, 12'hE49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE4C} : s_CHIP_23B_45132_reg = 8'h93;
         {3'b111, 12'hE4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE50} : s_CHIP_23B_45132_reg = 8'h94;
         {3'b111, 12'hE51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE54} : s_CHIP_23B_45132_reg = 8'h95;
         {3'b111, 12'hE55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE58} : s_CHIP_23B_45132_reg = 8'h96;
         {3'b111, 12'hE59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE5C} : s_CHIP_23B_45132_reg = 8'h97;
         {3'b111, 12'hE5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE60} : s_CHIP_23B_45132_reg = 8'h98;
         {3'b111, 12'hE61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE64} : s_CHIP_23B_45132_reg = 8'h99;
         {3'b111, 12'hE65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE68} : s_CHIP_23B_45132_reg = 8'h9A;
         {3'b111, 12'hE69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE6C} : s_CHIP_23B_45132_reg = 8'h9B;
         {3'b111, 12'hE6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE70} : s_CHIP_23B_45132_reg = 8'h9C;
         {3'b111, 12'hE71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE74} : s_CHIP_23B_45132_reg = 8'h9D;
         {3'b111, 12'hE75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE78} : s_CHIP_23B_45132_reg = 8'h9E;
         {3'b111, 12'hE79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE7C} : s_CHIP_23B_45132_reg = 8'h9F;
         {3'b111, 12'hE7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE80} : s_CHIP_23B_45132_reg = 8'hA0;
         {3'b111, 12'hE81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE84} : s_CHIP_23B_45132_reg = 8'hA1;
         {3'b111, 12'hE85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE88} : s_CHIP_23B_45132_reg = 8'hA2;
         {3'b111, 12'hE89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE8C} : s_CHIP_23B_45132_reg = 8'hA3;
         {3'b111, 12'hE8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE90} : s_CHIP_23B_45132_reg = 8'hA4;
         {3'b111, 12'hE91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE94} : s_CHIP_23B_45132_reg = 8'hA5;
         {3'b111, 12'hE95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE98} : s_CHIP_23B_45132_reg = 8'hA6;
         {3'b111, 12'hE99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hE9C} : s_CHIP_23B_45132_reg = 8'hA7;
         {3'b111, 12'hE9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEA0} : s_CHIP_23B_45132_reg = 8'hA8;
         {3'b111, 12'hEA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEA4} : s_CHIP_23B_45132_reg = 8'hA9;
         {3'b111, 12'hEA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEA8} : s_CHIP_23B_45132_reg = 8'hAA;
         {3'b111, 12'hEA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEAC} : s_CHIP_23B_45132_reg = 8'hAB;
         {3'b111, 12'hEAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEB0} : s_CHIP_23B_45132_reg = 8'hAC;
         {3'b111, 12'hEB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEB4} : s_CHIP_23B_45132_reg = 8'hAD;
         {3'b111, 12'hEB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEB8} : s_CHIP_23B_45132_reg = 8'hAE;
         {3'b111, 12'hEB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEBC} : s_CHIP_23B_45132_reg = 8'hAF;
         {3'b111, 12'hEBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEC0} : s_CHIP_23B_45132_reg = 8'hB0;
         {3'b111, 12'hEC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEC4} : s_CHIP_23B_45132_reg = 8'hB1;
         {3'b111, 12'hEC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEC8} : s_CHIP_23B_45132_reg = 8'hB2;
         {3'b111, 12'hEC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hECC} : s_CHIP_23B_45132_reg = 8'hB3;
         {3'b111, 12'hECD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hED0} : s_CHIP_23B_45132_reg = 8'hB4;
         {3'b111, 12'hED1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hED4} : s_CHIP_23B_45132_reg = 8'hB5;
         {3'b111, 12'hED5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hED8} : s_CHIP_23B_45132_reg = 8'hB6;
         {3'b111, 12'hED9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEDC} : s_CHIP_23B_45132_reg = 8'hB7;
         {3'b111, 12'hEDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEE0} : s_CHIP_23B_45132_reg = 8'hB8;
         {3'b111, 12'hEE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEE4} : s_CHIP_23B_45132_reg = 8'hB9;
         {3'b111, 12'hEE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEE8} : s_CHIP_23B_45132_reg = 8'hBA;
         {3'b111, 12'hEE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEEC} : s_CHIP_23B_45132_reg = 8'hBB;
         {3'b111, 12'hEED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEF0} : s_CHIP_23B_45132_reg = 8'hBC;
         {3'b111, 12'hEF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEF4} : s_CHIP_23B_45132_reg = 8'hBD;
         {3'b111, 12'hEF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEF8} : s_CHIP_23B_45132_reg = 8'hBE;
         {3'b111, 12'hEF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hEFC} : s_CHIP_23B_45132_reg = 8'hBF;
         {3'b111, 12'hEFD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF00} : s_CHIP_23B_45132_reg = 8'hC0;
         {3'b111, 12'hF01} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF04} : s_CHIP_23B_45132_reg = 8'hC1;
         {3'b111, 12'hF05} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF08} : s_CHIP_23B_45132_reg = 8'hC2;
         {3'b111, 12'hF09} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF0C} : s_CHIP_23B_45132_reg = 8'hC3;
         {3'b111, 12'hF0D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF10} : s_CHIP_23B_45132_reg = 8'hC4;
         {3'b111, 12'hF11} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF14} : s_CHIP_23B_45132_reg = 8'hC5;
         {3'b111, 12'hF15} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF18} : s_CHIP_23B_45132_reg = 8'hC6;
         {3'b111, 12'hF19} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF1C} : s_CHIP_23B_45132_reg = 8'hC7;
         {3'b111, 12'hF1D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF20} : s_CHIP_23B_45132_reg = 8'hC8;
         {3'b111, 12'hF21} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF24} : s_CHIP_23B_45132_reg = 8'hC9;
         {3'b111, 12'hF25} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF28} : s_CHIP_23B_45132_reg = 8'hCA;
         {3'b111, 12'hF29} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF2C} : s_CHIP_23B_45132_reg = 8'hCB;
         {3'b111, 12'hF2D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF30} : s_CHIP_23B_45132_reg = 8'hCC;
         {3'b111, 12'hF31} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF34} : s_CHIP_23B_45132_reg = 8'hCD;
         {3'b111, 12'hF35} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF38} : s_CHIP_23B_45132_reg = 8'hCE;
         {3'b111, 12'hF39} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF3C} : s_CHIP_23B_45132_reg = 8'hCF;
         {3'b111, 12'hF3D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF40} : s_CHIP_23B_45132_reg = 8'hD0;
         {3'b111, 12'hF41} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF44} : s_CHIP_23B_45132_reg = 8'hD1;
         {3'b111, 12'hF45} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF48} : s_CHIP_23B_45132_reg = 8'hD2;
         {3'b111, 12'hF49} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF4C} : s_CHIP_23B_45132_reg = 8'hD3;
         {3'b111, 12'hF4D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF50} : s_CHIP_23B_45132_reg = 8'hD4;
         {3'b111, 12'hF51} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF54} : s_CHIP_23B_45132_reg = 8'hD5;
         {3'b111, 12'hF55} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF58} : s_CHIP_23B_45132_reg = 8'hD6;
         {3'b111, 12'hF59} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF5C} : s_CHIP_23B_45132_reg = 8'hD7;
         {3'b111, 12'hF5D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF60} : s_CHIP_23B_45132_reg = 8'hD8;
         {3'b111, 12'hF61} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF64} : s_CHIP_23B_45132_reg = 8'hD9;
         {3'b111, 12'hF65} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF68} : s_CHIP_23B_45132_reg = 8'hDA;
         {3'b111, 12'hF69} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF6C} : s_CHIP_23B_45132_reg = 8'hDB;
         {3'b111, 12'hF6D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF70} : s_CHIP_23B_45132_reg = 8'hDC;
         {3'b111, 12'hF71} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF74} : s_CHIP_23B_45132_reg = 8'hDD;
         {3'b111, 12'hF75} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF78} : s_CHIP_23B_45132_reg = 8'hDE;
         {3'b111, 12'hF79} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF7C} : s_CHIP_23B_45132_reg = 8'hDF;
         {3'b111, 12'hF7D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF80} : s_CHIP_23B_45132_reg = 8'hE0;
         {3'b111, 12'hF81} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF84} : s_CHIP_23B_45132_reg = 8'hE1;
         {3'b111, 12'hF85} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF88} : s_CHIP_23B_45132_reg = 8'hE2;
         {3'b111, 12'hF89} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF8C} : s_CHIP_23B_45132_reg = 8'hE3;
         {3'b111, 12'hF8D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF90} : s_CHIP_23B_45132_reg = 8'hE4;
         {3'b111, 12'hF91} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF94} : s_CHIP_23B_45132_reg = 8'hE5;
         {3'b111, 12'hF95} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF98} : s_CHIP_23B_45132_reg = 8'hE6;
         {3'b111, 12'hF99} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hF9C} : s_CHIP_23B_45132_reg = 8'hE7;
         {3'b111, 12'hF9D} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFA0} : s_CHIP_23B_45132_reg = 8'hE8;
         {3'b111, 12'hFA1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFA4} : s_CHIP_23B_45132_reg = 8'hE9;
         {3'b111, 12'hFA5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFA8} : s_CHIP_23B_45132_reg = 8'hEA;
         {3'b111, 12'hFA9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFAC} : s_CHIP_23B_45132_reg = 8'hEB;
         {3'b111, 12'hFAD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFB0} : s_CHIP_23B_45132_reg = 8'hEC;
         {3'b111, 12'hFB1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFB4} : s_CHIP_23B_45132_reg = 8'hED;
         {3'b111, 12'hFB5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFB8} : s_CHIP_23B_45132_reg = 8'hEE;
         {3'b111, 12'hFB9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFBC} : s_CHIP_23B_45132_reg = 8'hEF;
         {3'b111, 12'hFBD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFC0} : s_CHIP_23B_45132_reg = 8'hF0;
         {3'b111, 12'hFC1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFC4} : s_CHIP_23B_45132_reg = 8'hF1;
         {3'b111, 12'hFC5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFC8} : s_CHIP_23B_45132_reg = 8'hF2;
         {3'b111, 12'hFC9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFCC} : s_CHIP_23B_45132_reg = 8'hF3;
         {3'b111, 12'hFCD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFD0} : s_CHIP_23B_45132_reg = 8'hF4;
         {3'b111, 12'hFD1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFD4} : s_CHIP_23B_45132_reg = 8'hF5;
         {3'b111, 12'hFD5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFD8} : s_CHIP_23B_45132_reg = 8'hF6;
         {3'b111, 12'hFD9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFDC} : s_CHIP_23B_45132_reg = 8'hF7;
         {3'b111, 12'hFDD} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFE0} : s_CHIP_23B_45132_reg = 8'hF8;
         {3'b111, 12'hFE1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFE4} : s_CHIP_23B_45132_reg = 8'hF9;
         {3'b111, 12'hFE5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFE8} : s_CHIP_23B_45132_reg = 8'hFA;
         {3'b111, 12'hFE9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFEC} : s_CHIP_23B_45132_reg = 8'hFB;
         {3'b111, 12'hFED} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFF0} : s_CHIP_23B_45132_reg = 8'hFC;
         {3'b111, 12'hFF1} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFF4} : s_CHIP_23B_45132_reg = 8'hFD;
         {3'b111, 12'hFF5} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFF8} : s_CHIP_23B_45132_reg = 8'hFE;
         {3'b111, 12'hFF9} : s_CHIP_23B_45132_reg = 8'h10;
         {3'b111, 12'hFFC} : s_CHIP_23B_45132_reg = 8'hFF;
         {3'b111, 12'hFFD} : s_CHIP_23B_45132_reg = 8'h10;
         default : s_CHIP_23B_45132_reg = 8'h00;
      endcase
   end

   assign s_databus[7:0] = s_CHIP_23B_45132_reg;

   // ROM: CHIP_26B_45133
   reg[7:0] s_CHIP_26B_45133_reg;
      always @(*)
      begin
         case (s_Address)
         {3'b000, 12'h000} : s_CHIP_26B_45133_reg = 8'hC4;
         {3'b000, 12'h003} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h004} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h007} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h008} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h00B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h00E} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h00F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h012} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h013} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h016} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h017} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h02B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h03A} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h03B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h03C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h03E} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'h03F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h040} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h041} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h043} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h045} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h047} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h048} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h049} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h04B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h04D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h04F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h051} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h052} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'h053} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h055} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h057} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h058} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h059} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h05B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h05E} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h05F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h060} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h061} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h062} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h063} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h065} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h067} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h069} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h06A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h06B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'h06D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h06F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h071} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h073} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h075} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h077} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'h079} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h07B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h07D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h07F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h081} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h083} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h084} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'h085} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h087} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h088} : s_CHIP_26B_45133_reg = 8'hC5;
         {3'b000, 12'h089} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h08B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h08C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b000, 12'h08D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h08F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h091} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h093} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h095} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h097} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h09B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'h09E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h09F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h0A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h0A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h0A8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h0A9} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h0AA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h0AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h0AC} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h0AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0AF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h0B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h0B5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h0B8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h0B9} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h0BA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h0BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h0BC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b000, 12'h0BD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h0BF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h0C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h0C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0C6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h0C7} : s_CHIP_26B_45133_reg = 8'hBB;
         {3'b000, 12'h0C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0CB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h0CC} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b000, 12'h0CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0CF} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b000, 12'h0D0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h0D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0D2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h0D3} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b000, 12'h0D4} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h0D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0D6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h0D7} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h0DB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h0DC} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'h0DF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h0E0} : s_CHIP_26B_45133_reg = 8'h58;
         {3'b000, 12'h0E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0E3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h0E4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b000, 12'h0E5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h0E7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h0E8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h0E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0EB} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b000, 12'h0EC} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h0ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h0EF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h0F0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h0F1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h0F2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h0F3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h0F7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'h104} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h105} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h106} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h107} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h108} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h109} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h10A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h10B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h10C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h10D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h10E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h10F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h110} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h111} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h112} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h113} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h115} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h116} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h117} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h119} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h11A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h11B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h11C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h11D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h11E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h11F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h120} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h121} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h122} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h123} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h125} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h126} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h127} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h129} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h12A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h12B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h12D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h12E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h12F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h131} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h132} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h133} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h135} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h136} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h137} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h139} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h13A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h13B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h13D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h13E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h13F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h141} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h142} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h143} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h145} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h146} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h147} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h149} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h14A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h14B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h14D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h14E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h14F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h151} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h152} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h153} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h155} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h156} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h157} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h159} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h15A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h15B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h15D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h15E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h15F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h161} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h162} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h163} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h165} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h166} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h167} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h169} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h16A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h16B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h16C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b000, 12'h16D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h16E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h16F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h170} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b000, 12'h171} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h172} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h173} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h174} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b000, 12'h175} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h176} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h177} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h178} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b000, 12'h179} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h17A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h17B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h17C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h17D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h17E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h17F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h180} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h181} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h182} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h183} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h184} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b000, 12'h185} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h186} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h187} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h188} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b000, 12'h189} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h18A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h18B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h18D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h18E} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b000, 12'h18F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h191} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h192} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h193} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h196} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h197} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h199} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h19B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h19C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h19D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h19F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h1A0} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h1A1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1A3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h1A4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h1A5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1A7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h1A8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'h1AA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1AB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h1AC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h1AD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1AF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h1B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h1B2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1B3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h1B6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1B7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h1B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h1BC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h1BE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1BF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h1C0} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h1C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1C3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h1C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1C7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h1C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h1CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h1CF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h1D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h1D2} : s_CHIP_26B_45133_reg = 8'h48;
         {3'b000, 12'h1D3} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'h1D4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h1D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h1D6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1D7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h1D8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h1D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h1DA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h1DB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h1DD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h1E2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1E3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h1E5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h1EA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1EB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h1ED} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h1F2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1F3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h1F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h1F8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h1FA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1FB} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'h1FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h1FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h200} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h202} : s_CHIP_26B_45133_reg = 8'h4C;
         {3'b000, 12'h203} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b000, 12'h205} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h207} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h208} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h20A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h20B} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'h20D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h20F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h210} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h212} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h213} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b000, 12'h215} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h217} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h218} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b000, 12'h219} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h21B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b000, 12'h21C} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b000, 12'h21D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h21F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h220} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b000, 12'h221} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h223} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h224} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b000, 12'h225} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h227} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h228} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b000, 12'h229} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h22B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h22D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h22E} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'h22F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h232} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h233} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h236} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h237} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b000, 12'h238} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h23B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h23C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h23F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h241} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h243} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h247} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h24B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h24E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h24F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h253} : s_CHIP_26B_45133_reg = 8'h7E;
         {3'b000, 12'h254} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h256} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h257} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'h259} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h25B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h25D} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b000, 12'h25E} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h25F} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b000, 12'h261} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h263} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h265} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b000, 12'h267} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h269} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h26B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h26D} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b000, 12'h26E} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h26F} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b000, 12'h271} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h273} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h275} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b000, 12'h276} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h277} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b000, 12'h278} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'h279} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h27B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'h27D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'h27E} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h27F} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b000, 12'h283} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h285} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h286} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h287} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h289} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h28B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h28D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h28F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h290} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h293} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h295} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'h297} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h299} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h29B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h29F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'h2A1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h2A3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h2A4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h2A7} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'h2A9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h2AB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h2AC} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h2AF} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b000, 12'h2B1} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h2B2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h2B3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h2B5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h2B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h2B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h2BB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h2BF} : s_CHIP_26B_45133_reg = 8'h1D;
         {3'b000, 12'h2C1} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h2C2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h2C3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h2C5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h2C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h2C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h2CB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h2CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h2CF} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b000, 12'h2D1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h2D3} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h2D5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h2D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h2DA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h2DB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h2DC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h2DD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h2DF} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h2E3} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h2E4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h2E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h2E7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h2E8} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h2E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h2EB} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'h2ED} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h2EF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h2F3} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b000, 12'h2F5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h2F6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h2F7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h2F9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h2FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h2FD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h2FF} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h300} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h301} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h303} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h305} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h307} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h308} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h309} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h30B} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'h30D} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h30E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h30F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h311} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h313} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h316} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h317} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h319} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h31A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h31B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h31D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h31F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h321} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h323} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h324} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h325} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h327} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h328} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h329} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h32B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h32C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h32F} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b000, 12'h331} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h332} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h333} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h335} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h337} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h33A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h33B} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h33D} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h33E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h33F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h341} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h343} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h345} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h347} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h348} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h349} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h34B} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h34C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h34D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h34F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h350} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h353} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b000, 12'h356} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h357} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'h359} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h35B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h35D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h35F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h361} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h363} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h365} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h367} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h369} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h36A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h36B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h36D} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h36F} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h371} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h372} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h373} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h375} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h377} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h378} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h379} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h37B} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b000, 12'h37D} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'h37F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h381} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'h383} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h384} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h385} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h387} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h389} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h38A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h38B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h38D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h38E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h38F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h391} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h392} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h393} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h395} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h396} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h397} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h399} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h39A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h39B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h39D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h39E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h39F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h3A3} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h3A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h3A6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h3A7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h3AA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h3AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3AD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3B1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3B2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h3B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3B4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3B5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h3B7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h3B8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h3B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h3BB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h3BD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h3BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h3BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3C1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3C5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3C9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3CD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3D1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3D5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3D9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3DD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h3DF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h3E1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h3E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3E5} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'h3E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3E9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'h3EB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h3EC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h3ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h3EF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h3F3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h3F5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h3F6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h3F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3F9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h3FC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h3FD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h3FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h402} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h403} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h405} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h407} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h409} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h40B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h40C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h40D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h40F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h411} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h413} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'h414} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h417} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b000, 12'h419} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h41B} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h41D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h41F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h421} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h423} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h425} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h427} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h429} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h42B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h42C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h42D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h42F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h432} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h433} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h434} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h435} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h437} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h439} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h43B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h43C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h43D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h43F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h440} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'h441} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h443} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h444} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h445} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h447} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h449} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h44B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h44C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h44D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h44F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'h450} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h451} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h453} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h455} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h457} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h459} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h45B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h45D} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'h45E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h45F} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h461} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h463} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h464} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'h465} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h467} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h469} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h46A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h46B} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b000, 12'h46C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h46D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h46F} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b000, 12'h471} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h472} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h473} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b000, 12'h475} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h476} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h477} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b000, 12'h478} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h479} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h47A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h47B} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b000, 12'h47C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h47D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h47F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h481} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h483} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b000, 12'h485} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h487} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h488} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h489} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h48B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h48D} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'h48E} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b000, 12'h48F} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b000, 12'h490} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h491} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'h492} : s_CHIP_26B_45133_reg = 8'hE8;
         {3'b000, 12'h493} : s_CHIP_26B_45133_reg = 8'hC4;
         {3'b000, 12'h495} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h497} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h498} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h499} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h49A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h49B} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'h49D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h49E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h49F} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h4A0} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h4A1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h4A3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h4A4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h4A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h4A7} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h4A8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h4A9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h4AB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h4AC} : s_CHIP_26B_45133_reg = 8'hD1;
         {3'b000, 12'h4AD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h4AF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h4B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h4B2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h4B3} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b000, 12'h4B4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h4B5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h4B7} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h4B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h4BA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h4BB} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b000, 12'h4BC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h4BD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h4BF} : s_CHIP_26B_45133_reg = 8'h38;
         {3'b000, 12'h4C1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h4C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h4C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h4C6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h4C7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h4C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h4CB} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b000, 12'h4CC} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h4CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h4CF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h4D1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h4D3} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'h4D4} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b000, 12'h4D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h4D7} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h4D8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h4D9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h4DB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h4DE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h4DF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h4E0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h4E2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h4E3} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'h4E5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h4E7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h4E8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h4E9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h4EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h4EE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h4EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h4F0} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h4F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h4F2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h4F3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h4F4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h4F5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h4F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h4FA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h4FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h4FC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h4FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h4FF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h500} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h501} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h503} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h504} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h505} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h506} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h507} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b000, 12'h509} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h50B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h50C} : s_CHIP_26B_45133_reg = 8'h91;
         {3'b000, 12'h50D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h50E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h50F} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b000, 12'h511} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h512} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h513} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h514} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h515} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h517} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h518} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h519} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h51B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h51C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h51D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h51E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h51F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h521} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h523} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h524} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b000, 12'h525} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h527} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h528} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b000, 12'h529} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h52B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h52C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h52D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h52F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h531} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h533} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h535} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h537} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h539} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h53B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h53D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h53E} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'h53F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h541} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h543} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b000, 12'h544} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h545} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h546} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h547} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h548} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b000, 12'h549} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h54A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h54B} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b000, 12'h54C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h54D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h54E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h54F} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b000, 12'h551} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h552} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h553} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h554} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h555} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'h556} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h557} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h559} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'h55A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h55B} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b000, 12'h55C} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'h55D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h55F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h561} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h562} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h563} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h564} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h565} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h567} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h568} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'h569} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h56B} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h56C} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b000, 12'h56D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h56F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h570} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h573} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h574} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h575} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h577} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h578} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h579} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h57B} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'h57C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'h57D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h57F} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h581} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'h583} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h584} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h585} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h587} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'h589} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h58B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h58C} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b000, 12'h58D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h58F} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h590} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'h591} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h593} : s_CHIP_26B_45133_reg = 8'h7E;
         {3'b000, 12'h595} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h596} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b000, 12'h597} : s_CHIP_26B_45133_reg = 8'hBB;
         {3'b000, 12'h599} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h59B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h59D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h59F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h5A0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h5A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5A3} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'h5A4} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b000, 12'h5A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5A7} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'h5A8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h5A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5AA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h5AB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'h5AC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h5AD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h5AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h5B0} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b000, 12'h5B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5B3} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'h5B4} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'h5B5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h5B6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h5B7} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h5B8} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'h5B9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h5BB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h5BC} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b000, 12'h5BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5BF} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'h5C0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h5C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h5C4} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h5C5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h5C7} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b000, 12'h5C8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h5C9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h5CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h5CC} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b000, 12'h5CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5CF} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'h5D0} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b000, 12'h5D1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h5D2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h5D3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h5D4} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h5D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5D7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h5D8} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h5D9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h5DA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h5DB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'h5DC} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b000, 12'h5DD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h5DE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h5DF} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b000, 12'h5E0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h5E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5E2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h5E3} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b000, 12'h5E4} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b000, 12'h5E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5E7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h5E8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'h5E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5EB} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h5ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5EF} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h5F0} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b000, 12'h5F3} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h5F5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h5F6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h5F7} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h5F8} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b000, 12'h5F9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h5FB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h5FC} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h5FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h5FF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h600} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h601} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h603} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h604} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h605} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'h607} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h608} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h609} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h60A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h60B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'h60C} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b000, 12'h60D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h60F} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b000, 12'h610} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h612} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h613} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b000, 12'h615} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h617} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h618} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h61B} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b000, 12'h61C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h61D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h61E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h61F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'h620} : s_CHIP_26B_45133_reg = 8'hD1;
         {3'b000, 12'h621} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h623} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h625} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h626} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h627} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b000, 12'h628} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h629} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h62B} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h62C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h62D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h62F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h630} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h632} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h633} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b000, 12'h635} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h637} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h638} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h639} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h63B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h63C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h63D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h63E} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'h63F} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b000, 12'h640} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h641} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h642} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'h643} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b000, 12'h644} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h645} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h647} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h64B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h64D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h64F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h650} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h651} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h653} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h654} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h655} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h656} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'h657} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b000, 12'h658} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h659} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h65A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'h65B} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b000, 12'h65C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h65D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h65F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h663} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h665} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h666} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h667} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h669} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h66A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'h66B} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b000, 12'h66C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h66D} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h66F} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b000, 12'h670} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h671} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h673} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h675} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h677} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h678} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h67B} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b000, 12'h67C} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b000, 12'h67D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h67F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h680} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h681} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h683} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h686} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h687} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h688} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b000, 12'h689} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h68B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h68C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h68D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h68F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h692} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h693} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h694} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h695} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h697} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b000, 12'h69B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h69C} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b000, 12'h69D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h69F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h6A0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h6A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6A4} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b000, 12'h6A5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h6A7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h6A8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h6AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6AC} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h6AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h6AE} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h6AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6B5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h6B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6BD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h6BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6C0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h6C1} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h6C3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h6C4} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'h6C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h6C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6C8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h6CB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h6CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h6CF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h6D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h6D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6D4} : s_CHIP_26B_45133_reg = 8'hF2;
         {3'b000, 12'h6D5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h6D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6DA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h6DB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h6DC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'h6DD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h6DF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h6E1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h6E2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h6E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6E6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h6E7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h6E8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'h6E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h6EB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h6EC} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h6ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h6EE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h6EF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h6F0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h6F1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h6F3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h6F5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h6F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6F8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h6F9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h6FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h6FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h6FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h703} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h704} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h705} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h707} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h708} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'h709} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h70A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h70B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h70C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h70D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h70E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h70F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b000, 12'h710} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h711} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h713} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h714} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h715} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h717} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h718} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h719} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h71B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h71C} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b000, 12'h71D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h71F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h720} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h721} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h723} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h725} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h726} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h727} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h728} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h729} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h72B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h72C} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b000, 12'h72D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h72F} : s_CHIP_26B_45133_reg = 8'h3D;
         {3'b000, 12'h730} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b000, 12'h731} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h733} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h735} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h737} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b000, 12'h738} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h739} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h73A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h73B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h73D} : s_CHIP_26B_45133_reg = 8'h95;
         {3'b000, 12'h73E} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'h73F} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b000, 12'h740} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h741} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h743} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b000, 12'h744} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h745} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h747} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h749} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h74B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h74C} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b000, 12'h74D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h74F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h750} : s_CHIP_26B_45133_reg = 8'hD1;
         {3'b000, 12'h753} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h754} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h755} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h756} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h757} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h758} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h759} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h75B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h75C} : s_CHIP_26B_45133_reg = 8'h3F;
         {3'b000, 12'h75D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h75F} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h760} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h761} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h763} : s_CHIP_26B_45133_reg = 8'h3D;
         {3'b000, 12'h765} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h767} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h768} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h769} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'h76A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h76B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h76C} : s_CHIP_26B_45133_reg = 8'h91;
         {3'b000, 12'h76D} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b000, 12'h76F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h770} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'h771} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h772} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h773} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'h775} : s_CHIP_26B_45133_reg = 8'h95;
         {3'b000, 12'h777} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b000, 12'h778} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h77B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b000, 12'h77D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h77E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h77F} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h780} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h781} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h783} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h785} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h787} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h788} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b000, 12'h789} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h78B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h78D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h78F} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h790} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b000, 12'h791} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h793} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h795} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h797} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h798} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h799} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h79B} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h79D} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h79E} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h79F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h7A0} : s_CHIP_26B_45133_reg = 8'hD7;
         {3'b000, 12'h7A1} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h7A3} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b000, 12'h7A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h7A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h7AC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h7AD} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'h7AE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h7AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h7B1} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h7B3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h7B4} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'h7B5} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h7B8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h7B9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h7BB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h7BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7BF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h7C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7C3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h7C4} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h7C5} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h7C7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h7C8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h7C9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h7CB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h7CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7CF} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h7D0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h7D1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h7D3} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b000, 12'h7D4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b000, 12'h7D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7D7} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h7D8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h7D9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h7DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h7DC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h7DE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h7DF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h7E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7E2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h7E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h7E4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h7E5} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'h7E7} : s_CHIP_26B_45133_reg = 8'hFA;
         {3'b000, 12'h7E9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'h7EB} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b000, 12'h7EC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'h7ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7EF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h7F1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h7F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h7F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7F7} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h7F8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h7F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h7FB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h7FD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h7FF} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h800} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h801} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b000, 12'h803} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'h804} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'h805} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h807} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h809} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h80B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h80C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h80D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h80F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h813} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h814} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'h815} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h817} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b000, 12'h818} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b000, 12'h819} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h81B} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h81C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'h81D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h81F} : s_CHIP_26B_45133_reg = 8'hEF;
         {3'b000, 12'h820} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h821} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h822} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h823} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h824} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h825} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h827} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h828} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h829} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h82B} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h82C} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b000, 12'h82D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h830} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h831} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h833} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h834} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h835} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h837} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h838} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h839} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h83B} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'h83C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h83D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h83F} : s_CHIP_26B_45133_reg = 8'h3D;
         {3'b000, 12'h840} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h841} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h843} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h844} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h845} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h846} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h847} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h849} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h84B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h84C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h84D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h84F} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'h850} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h851} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h853} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'h854} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h855} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h857} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h858} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h859} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h85B} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'h85C} : s_CHIP_26B_45133_reg = 8'hE2;
         {3'b000, 12'h85F} : s_CHIP_26B_45133_reg = 8'h3D;
         {3'b000, 12'h860} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h861} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h862} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h863} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h864} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'h865} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h867} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h868} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h869} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h86B} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b000, 12'h86C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h86F} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h870} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'h871} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h873} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h875} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h876} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h877} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h878} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h879} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h87B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h87D} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h87E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'h87F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h880} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h881} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h883} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b000, 12'h884} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h885} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h886} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h887} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h888} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h889} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h88B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h88C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h88D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h88F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h891} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h893} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h895} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h896} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b000, 12'h897} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h899} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h89A} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b000, 12'h89B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h89C} : s_CHIP_26B_45133_reg = 8'h3F;
         {3'b000, 12'h89D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h89F} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h8A0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h8A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h8A3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h8A4} : s_CHIP_26B_45133_reg = 8'hA2;
         {3'b000, 12'h8A7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h8A8} : s_CHIP_26B_45133_reg = 8'h3F;
         {3'b000, 12'h8A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h8AB} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h8AC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h8AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h8AF} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h8B0} : s_CHIP_26B_45133_reg = 8'hA2;
         {3'b000, 12'h8B3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h8B4} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'h8B5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h8B6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h8B7} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b000, 12'h8B8} : s_CHIP_26B_45133_reg = 8'hF2;
         {3'b000, 12'h8B9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h8BB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h8BC} : s_CHIP_26B_45133_reg = 8'hE2;
         {3'b000, 12'h8BD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h8BF} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b000, 12'h8C1} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h8C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h8C4} : s_CHIP_26B_45133_reg = 8'hB2;
         {3'b000, 12'h8C5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h8C7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h8C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h8CB} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h8CC} : s_CHIP_26B_45133_reg = 8'hB2;
         {3'b000, 12'h8CD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h8CF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h8D0} : s_CHIP_26B_45133_reg = 8'h3F;
         {3'b000, 12'h8D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h8D3} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h8D4} : s_CHIP_26B_45133_reg = 8'hF2;
         {3'b000, 12'h8D5} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b000, 12'h8D6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h8D7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'h8D8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h8D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h8DB} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b000, 12'h8DC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'h8DD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h8DF} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b000, 12'h8E0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h8E1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h8E3} : s_CHIP_26B_45133_reg = 8'h38;
         {3'b000, 12'h8E4} : s_CHIP_26B_45133_reg = 8'hE2;
         {3'b000, 12'h8E5} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'h8E6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h8E7} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'h8E9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h8EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h8ED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h8EF} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h8F0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h8F1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h8F2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h8F3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h8F4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h8F5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h8F6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h8F7} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'h8FA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h8FB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h8FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h8FF} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'h900} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h901} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h903} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h905} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h907} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b000, 12'h908} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h909} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h90A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'h90B} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b000, 12'h90C} : s_CHIP_26B_45133_reg = 8'hF2;
         {3'b000, 12'h90D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h90F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h910} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h911} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h912} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'h913} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b000, 12'h914} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h915} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h917} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h919} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h91A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'h91B} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b000, 12'h91C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h91D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h91F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h920} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h921} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h923} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h924} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h925} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h927} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h929} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h92B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h92C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'h92D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h92E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h92F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h930} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h931} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h933} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h935} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b000, 12'h937} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b000, 12'h938} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h939} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b000, 12'h93B} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b000, 12'h93C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h93D} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'h93F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h941} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'h943} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b000, 12'h944} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h946} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h947} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h948} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h949} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h94B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h94C} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b000, 12'h94F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h951} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h953} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'h954} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'h955} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h957} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h959} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h95B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h95C} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b000, 12'h95D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h95F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h962} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h963} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h964} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h965} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h967} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'h96A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h96B} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b000, 12'h96D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h96F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h970} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h971} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h972} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h973} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h975} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h977} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h978} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h979} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h97B} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b000, 12'h97C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h97D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h97F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h981} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h983} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h985} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h987} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h988} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'h989} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h98B} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h98D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h98F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h990} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h991} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h992} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'h993} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h994} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h995} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h997} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h998} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'h999} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h99B} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b000, 12'h99D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h99F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h9A1} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'h9A3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h9A5} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'h9A7} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b000, 12'h9A8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'h9A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9AB} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b000, 12'h9AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9AF} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b000, 12'h9B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h9B4} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'h9B5} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'h9B7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h9B9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'h9BB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h9BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9BE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'h9BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h9C1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h9C3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'h9C4} : s_CHIP_26B_45133_reg = 8'h3F;
         {3'b000, 12'h9C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9C7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h9C8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h9C9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h9CB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h9CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9CF} : s_CHIP_26B_45133_reg = 8'hB3;
         {3'b000, 12'h9D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'h9D1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h9D3} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h9D4} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'h9D5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h9D7} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'h9D9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'h9DB} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b000, 12'h9DD} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'h9DE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'h9DF} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b000, 12'h9E0} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b000, 12'h9E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9E3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'h9E5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h9E7} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'h9E8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'h9E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9EB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'h9ED} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'h9EE} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b000, 12'h9EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h9F0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'h9F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9F2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'h9F3} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'h9F5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'h9F7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'h9F8} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h9F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'h9FB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'h9FC} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'h9FD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'h9FF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hA01} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA02} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA03} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hA05} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA07} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hA08} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hA09} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hA0B} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b000, 12'hA0D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA0F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hA11} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA12} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA13} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hA15} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA17} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hA19} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA1B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hA1D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hA1F} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'hA20} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b000, 12'hA21} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hA22} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA23} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'hA24} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hA25} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hA26} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA27} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hA29} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA2B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hA2C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hA2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA2E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA2F} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'hA30} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hA31} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA32} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hA33} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hA34} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hA35} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hA37} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hA38} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b000, 12'hA39} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA3A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA3B} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'hA3D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA3E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hA3F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hA40} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hA41} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hA43} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hA44} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hA45} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hA46} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA47} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'hA48} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hA49} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA4A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA4B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hA4C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hA4D} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hA4E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA4F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hA51} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA53} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'hA55} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA56} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b000, 12'hA57} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b000, 12'hA58} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hA59} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA5B} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b000, 12'hA5C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'hA5D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA5E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA5F} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'hA60} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hA61} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA63} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hA65} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA67} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hA69} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA6B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hA6C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA6E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA6F} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'hA71} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA72} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hA73} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'hA74} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'hA75} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hA77} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b000, 12'hA78} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA79} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA7A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA7B} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'hA7C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hA7D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA7E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hA7F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hA80} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hA81} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA82} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA83} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b000, 12'hA84} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA85} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA86} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA87} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'hA88} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA89} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'hA8A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hA8B} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hA8D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA8F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hA90} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hA91} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA92} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA93} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'hA94} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hA95} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hA96} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hA97} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hA98} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hA99} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA9B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hA9C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hA9D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hA9E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hA9F} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'hAA1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hAA2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hAA3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hAA5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAA7} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b000, 12'hAA9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAAB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'hAAD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hAAE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hAAF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'hAB1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAB3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hAB4} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hAB5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAB6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hAB7} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b000, 12'hAB9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hABA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hABB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hABD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hABF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hAC0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'hAC1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAC3} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b000, 12'hAC5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hAC6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hAC7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hAC8} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hAC9} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hACB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hACC} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hACE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'hACF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hAD0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'hAD1} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'hAD3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hAD4} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hAD5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAD7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hAD8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'hAD9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hADB} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hADC} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'hADD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hADF} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b000, 12'hAE0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'hAE1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAE3} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hAE4} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hAE5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAE7} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hAE8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'hAE9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hAEA} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAEB} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hAEC} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hAED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hAEF} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hAF0} : s_CHIP_26B_45133_reg = 8'hB2;
         {3'b000, 12'hAF1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hAF3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hAF4} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hAF5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hAF6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hAF7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hAF9} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'hAFB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hAFC} : s_CHIP_26B_45133_reg = 8'h82;
         {3'b000, 12'hAFD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hAFF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hB00} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hB01} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hB03} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hB04} : s_CHIP_26B_45133_reg = 8'hB2;
         {3'b000, 12'hB05} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hB07} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hB09} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hB0A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hB0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hB0D} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hB0F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hB10} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hB11} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hB13} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hB14} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hB15} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hB16} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hB17} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hB18} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'hB19} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hB1B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hB1C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hB1D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB1F} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'hB20} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hB21} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hB23} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hB24} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hB27} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hB28} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hB29} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hB2A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hB2B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hB2C} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'hB2D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hB2F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hB30} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hB31} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB33} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'hB34} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hB35} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hB37} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hB38} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hB3B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hB3C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hB3D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hB3F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hB41} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB43} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hB44} : s_CHIP_26B_45133_reg = 8'h82;
         {3'b000, 12'hB45} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hB47} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hB49} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB4B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hB4D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB4F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hB51} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hB53} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hB54} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hB55} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hB57} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hB59} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB5B} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b000, 12'hB5C} : s_CHIP_26B_45133_reg = 8'h82;
         {3'b000, 12'hB5D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hB5F} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hB60} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hB61} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB62} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hB63} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hB64} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hB65} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB67} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b000, 12'hB68} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hB6A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hB6B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hB6C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'hB6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB6F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hB70} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b000, 12'hB71} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB73} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hB74} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hB75} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hB77} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hB78} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'hB79} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hB7B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hB7C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hB7D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hB7E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hB7F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hB80} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hB81} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hB83} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b000, 12'hB84} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'hB85} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB87} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hB88} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b000, 12'hB89} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hB8A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hB8B} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hB8C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hB8D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB8F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hB90} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hB91} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB93} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hB94} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'hB95} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB97} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hB9A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hB9B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hB9D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hB9F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hBA1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBA3} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hBA5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hBA6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hBA7} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b000, 12'hBA8} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b000, 12'hBA9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hBAB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hBAC} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b000, 12'hBAD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hBAF} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hBB0} : s_CHIP_26B_45133_reg = 8'hA2;
         {3'b000, 12'hBB1} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'hBB3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hBB4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hBB5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hBB6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hBB7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hBB9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hBBB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hBBC} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b000, 12'hBBF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hBC0} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hBC1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBC2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hBC3} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'hBC4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hBC5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBC6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hBC7} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hBC8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hBC9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBCA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hBCB} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b000, 12'hBCC} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hBCD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBCF} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'hBD0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hBD1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBD2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hBD3} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b000, 12'hBD4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'hBD5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBD7} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hBDB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hBDC} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hBDD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hBDF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hBE1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBE2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hBE3} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'hBE5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBE7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hBE8} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hBEB} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b000, 12'hBED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBEF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hBF0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hBF1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hBF3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hBF4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hBF7} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b000, 12'hBF8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hBF9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hBFB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hBFD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hBFE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hBFF} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b000, 12'hC01} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC03} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hC04} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hC07} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b000, 12'hC08} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hC09} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hC0C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hC0F} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hC10} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hC11} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC13} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hC14} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hC15} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hC17} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC18} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hC19} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hC1B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hC1C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hC1F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hC20} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hC21} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC23} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hC24} : s_CHIP_26B_45133_reg = 8'hC3;
         {3'b000, 12'hC27} : s_CHIP_26B_45133_reg = 8'h77;
         {3'b000, 12'hC28} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hC29} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC2B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hC2C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hC2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC2F} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hC30} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b000, 12'hC31} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC33} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hC34} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hC35} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hC37} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hC38} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hC39} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC3B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hC3C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hC3D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC3F} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC40} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b000, 12'hC41} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hC43} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hC44} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hC45} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC47} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hC48} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hC49} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC4B} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC4C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hC4D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hC4F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hC50} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hC51} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hC52} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hC53} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b000, 12'hC54} : s_CHIP_26B_45133_reg = 8'hC3;
         {3'b000, 12'hC55} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hC57} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b000, 12'hC58} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'hC59} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC5B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hC5C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hC5D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hC5F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hC60} : s_CHIP_26B_45133_reg = 8'h93;
         {3'b000, 12'hC61} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hC63} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hC64} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hC65} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC67} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hC68} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hC69} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC6B} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hC6C} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hC6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC6F} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hC70} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hC71} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC73} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hC74} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC75} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC77} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b000, 12'hC78} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hC79} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hC7B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hC7C} : s_CHIP_26B_45133_reg = 8'hE3;
         {3'b000, 12'hC7D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hC7F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hC81} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hC82} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hC83} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'hC84} : s_CHIP_26B_45133_reg = 8'h52;
         {3'b000, 12'hC85} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC87} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'hC88} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'hC89} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC8B} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'hC8C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hC8D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC8E} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hC8F} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'hC90} : s_CHIP_26B_45133_reg = 8'h53;
         {3'b000, 12'hC91} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC93} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'hC94} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'hC95} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC97} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b000, 12'hC98} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hC99} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC9B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hC9C} : s_CHIP_26B_45133_reg = 8'h53;
         {3'b000, 12'hC9D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hC9F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hCA0} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'hCA1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hCA3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hCA4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hCA5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hCA7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hCA8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hCA9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hCAB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hCAC} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b000, 12'hCAD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hCAF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hCB0} : s_CHIP_26B_45133_reg = 8'hD3;
         {3'b000, 12'hCB1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hCB3} : s_CHIP_26B_45133_reg = 8'hA6;
         {3'b000, 12'hCB4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hCB5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hCB6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hCB7} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'hCB8} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b000, 12'hCB9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hCBB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hCBC} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b000, 12'hCBD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hCBF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hCC1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hCC2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hCC3} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hCC5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hCC6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hCC7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hCC8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hCC9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hCCB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hCCC} : s_CHIP_26B_45133_reg = 8'h93;
         {3'b000, 12'hCCD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hCCF} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b000, 12'hCD0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hCD3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hCD4} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'hCD5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hCD7} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b000, 12'hCD8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hCD9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'hCDB} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hCDC} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hCDD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hCDF} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hCE0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hCE1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hCE2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hCE3} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hCE4} : s_CHIP_26B_45133_reg = 8'h82;
         {3'b000, 12'hCE5} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b000, 12'hCE7} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hCE8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hCE9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hCEB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hCEC} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hCED} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hCEE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hCEF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hCF0} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b000, 12'hCF1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hCF3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hCF5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hCF7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hCF8} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hCFB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hCFC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hCFD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hCFE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hCFF} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b000, 12'hD00} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b000, 12'hD01} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hD03} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hD04} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD05} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD07} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hD08} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hD0C} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'hD0D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD0F} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b000, 12'hD10} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hD11} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'hD13} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hD14} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hD15} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hD17} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hD18} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hD19} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hD1A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hD1B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hD1C} : s_CHIP_26B_45133_reg = 8'hC3;
         {3'b000, 12'hD1D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hD1F} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hD20} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hD21} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD23} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hD24} : s_CHIP_26B_45133_reg = 8'hC3;
         {3'b000, 12'hD25} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD27} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hD28} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD2B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hD2C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD2D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD2F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hD30} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD31} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD33} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hD36} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hD37} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hD38} : s_CHIP_26B_45133_reg = 8'hD3;
         {3'b000, 12'hD39} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hD3B} : s_CHIP_26B_45133_reg = 8'hA6;
         {3'b000, 12'hD3C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hD3D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hD3E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hD3F} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b000, 12'hD40} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b000, 12'hD41} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b000, 12'hD43} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hD44} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b000, 12'hD45} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD47} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b000, 12'hD48} : s_CHIP_26B_45133_reg = 8'h93;
         {3'b000, 12'hD49} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD4B} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hD4C} : s_CHIP_26B_45133_reg = 8'hC3;
         {3'b000, 12'hD4D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD4F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hD50} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD51} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD53} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'hD54} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hD55} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hD56} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hD57} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hD58} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b000, 12'hD59} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hD5B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hD5E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hD5F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hD60} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'hD61} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD63} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b000, 12'hD64} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hD65} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'hD67} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hD68} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hD69} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hD6B} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hD6C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hD6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hD6E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hD6F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hD70} : s_CHIP_26B_45133_reg = 8'h83;
         {3'b000, 12'hD71} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hD73} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hD74} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD75} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD77} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hD78} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD79} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD7B} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b000, 12'hD7C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hD7D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hD7F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hD80} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b000, 12'hD81} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD83} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hD84} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD86} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hD87} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hD88} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hD89} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD8B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hD8C} : s_CHIP_26B_45133_reg = 8'hC3;
         {3'b000, 12'hD8D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD8F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hD90} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD93} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hD94} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hD95} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hD96} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hD97} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b000, 12'hD98} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b000, 12'hD99} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b000, 12'hD9B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hD9C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hD9D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hD9F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hDA0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hDA1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hDA3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hDA4} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hDA5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hDA6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hDA7} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hDA8} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hDA9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hDAB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hDAE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hDAF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hDB0} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b000, 12'hDB1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hDB3} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b000, 12'hDB5} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'hDB7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hDB8} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hDB9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hDBB} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hDBC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hDBD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDBE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hDBF} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hDC0} : s_CHIP_26B_45133_reg = 8'hC2;
         {3'b000, 12'hDC1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hDC3} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hDC4} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hDC5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hDC7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hDC8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hDC9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hDCB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hDCE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hDCF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hDD0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'hDD1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hDD3} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'hDD4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hDD5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hDD7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hDD8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hDD9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDDB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hDDC} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'hDDD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hDDF} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b000, 12'hDE0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hDE1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDE2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hDE3} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b000, 12'hDE4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hDE5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDE7} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b000, 12'hDE8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hDE9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDEC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'hDED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDEF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hDF0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hDF1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDF3} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'hDF4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hDF5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDF6} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDF7} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hDF8} : s_CHIP_26B_45133_reg = 8'hB3;
         {3'b000, 12'hDF9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hDFB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hDFD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hDFE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hDFF} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b000, 12'hE01} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'hE02} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hE03} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hE04} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hE05} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hE06} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE07} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b000, 12'hE08} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hE09} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b000, 12'hE0B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'hE0C} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b000, 12'hE0D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hE0F} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'hE10} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE11} : s_CHIP_26B_45133_reg = 8'h91;
         {3'b000, 12'hE13} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hE14} : s_CHIP_26B_45133_reg = 8'hC3;
         {3'b000, 12'hE15} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hE16} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hE17} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b000, 12'hE18} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hE19} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE1B} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b000, 12'hE1D} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'hE1F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b000, 12'hE20} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE21} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b000, 12'hE23} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hE24} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hE25} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'hE27} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hE28} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hE29} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE2A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE2B} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'hE2C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hE2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE2E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE2F} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE30} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hE31} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE32} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE33} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b000, 12'hE34} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE35} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hE37} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b000, 12'hE38} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b000, 12'hE39} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hE3A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE3B} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE3C} : s_CHIP_26B_45133_reg = 8'h93;
         {3'b000, 12'hE3E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE3F} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b000, 12'hE40} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hE41} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE42} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE43} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'hE45} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE46} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE47} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b000, 12'hE48} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'hE49} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE4A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE4B} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b000, 12'hE4F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hE50} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hE51} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE53} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hE54} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE57} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b000, 12'hE58} : s_CHIP_26B_45133_reg = 8'hD3;
         {3'b000, 12'hE59} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hE5A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hE5B} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hE5C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE5D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hE5F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hE60} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hE61} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE63} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'hE64} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hE65} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hE67} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hE68} : s_CHIP_26B_45133_reg = 8'hCF;
         {3'b000, 12'hE69} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE6B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hE6C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE6F} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hE70} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hE71} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE72} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE73} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b000, 12'hE74} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b000, 12'hE75} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hE76} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hE77} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b000, 12'hE78} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b000, 12'hE79} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE7B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hE7C} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b000, 12'hE7D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hE7E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hE7F} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'hE80} : s_CHIP_26B_45133_reg = 8'hCF;
         {3'b000, 12'hE81} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE83} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hE84} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE85} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE87} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hE88} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hE89} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE8B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hE8C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hE8D} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hE8F} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hE90} : s_CHIP_26B_45133_reg = 8'hB2;
         {3'b000, 12'hE91} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hE93} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hE94} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hE95} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE97} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE98} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b000, 12'hE99} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE9A} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE9B} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hE9C} : s_CHIP_26B_45133_reg = 8'hEF;
         {3'b000, 12'hE9D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hE9F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hEA0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hEA1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hEA3} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hEA4} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b000, 12'hEA5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hEA7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hEA8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hEA9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hEAB} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hEAC} : s_CHIP_26B_45133_reg = 8'hA3;
         {3'b000, 12'hEAD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hEAF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hEB1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hEB2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hEB3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hEB5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hEB7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hEB8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hEB9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hEBB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hEBD} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'hEBE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hEBF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hEC1} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'hEC3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hEC4} : s_CHIP_26B_45133_reg = 8'hD3;
         {3'b000, 12'hEC5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hEC7} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hEC8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hEC9} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'hECB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hECC} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hECD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hECF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hED0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hED1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hED2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hED3} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hED5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hED6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hED7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hED8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hEDB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hEDC} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b000, 12'hEDD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hEDF} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hEE0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hEE1} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'hEE3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hEE4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hEE5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hEE7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hEE8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hEE9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hEEB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hEED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hEEF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hEF0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hEF3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hEF4} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hEF5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hEF7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hEF9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hEFB} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hEFD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hEFE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hEFF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b000, 12'hF01} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF02} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hF03} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hF04} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b000, 12'hF05} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hF07} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hF08} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF09} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'hF0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hF0D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF0E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hF0F} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'hF11} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF13} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hF14} : s_CHIP_26B_45133_reg = 8'h82;
         {3'b000, 12'hF15} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hF17} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hF18} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF19} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hF1B} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b000, 12'hF1C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF1D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hF1E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hF1F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b000, 12'hF20} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF23} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hF24} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF25} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hF27} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hF28} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF29} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF2B} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b000, 12'hF2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF2E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hF2F} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b000, 12'hF30} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b000, 12'hF31} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hF33} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b000, 12'hF34} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF35} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'hF37} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hF39} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF3A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hF3B} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b000, 12'hF3D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF3F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hF41} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF43} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b000, 12'hF44} : s_CHIP_26B_45133_reg = 8'h82;
         {3'b000, 12'hF45} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hF47} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b000, 12'hF48} : s_CHIP_26B_45133_reg = 8'hE3;
         {3'b000, 12'hF49} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hF4B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hF4C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF4D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hF4F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hF50} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF53} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hF54} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'hF55} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hF56} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hF57} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hF59} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF5A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hF5B} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b000, 12'hF5C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'hF5D} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b000, 12'hF5F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b000, 12'hF61} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'hF63} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hF64} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF65} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b000, 12'hF67} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'hF69} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b000, 12'hF6B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hF6D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'hF6F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hF70} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hF71} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b000, 12'hF73} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hF74} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b000, 12'hF75} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hF76} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b000, 12'hF77} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b000, 12'hF78} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b000, 12'hF79} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b000, 12'hF7A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hF7B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hF7C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF7D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hF7F} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'hF81} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'hF82} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'hF83} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hF85} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF87} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hF89} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hF8A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hF8B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hF8C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF8D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b000, 12'hF8F} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'hF91} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b000, 12'hF92} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'hF93} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b000, 12'hF95} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hF96} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hF97} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b000, 12'hF99} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hF9B} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hF9C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hF9D} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'hF9F} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hFA0} : s_CHIP_26B_45133_reg = 8'hA3;
         {3'b000, 12'hFA1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hFA3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hFA4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hFA5} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b000, 12'hFA6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hFA7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hFA8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hFA9} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b000, 12'hFAB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hFAC} : s_CHIP_26B_45133_reg = 8'hB3;
         {3'b000, 12'hFAD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hFAF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hFB0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hFB1} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b000, 12'hFB2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hFB3} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b000, 12'hFB4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hFB5} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b000, 12'hFB7} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b000, 12'hFB8} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b000, 12'hFB9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hFBB} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b000, 12'hFBC} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b000, 12'hFBD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hFBF} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b000, 12'hFC1} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b000, 12'hFC3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hFC5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b000, 12'hFC7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b000, 12'hFC8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b000, 12'hFC9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b000, 12'hFCA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b000, 12'hFCB} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hFCD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hFCF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hFD0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b000, 12'hFD1} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b000, 12'hFD3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b000, 12'hFD6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'hFD7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hFDA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'hFDB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hFDD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hFDF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hFE1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hFE2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hFE3} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b000, 12'hFE5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hFE6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'hFE7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b000, 12'hFEA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'hFEB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b000, 12'hFED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hFEE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b000, 12'hFEF} : s_CHIP_26B_45133_reg = 8'hFB;
         {3'b000, 12'hFF0} : s_CHIP_26B_45133_reg = 8'hFE;
         {3'b000, 12'hFF2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'hFF3} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b000, 12'hFF5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b000, 12'hFF6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hFF7} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b000, 12'hFF8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b000, 12'hFF9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b000, 12'hFFA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b000, 12'hFFB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b000, 12'hFFC} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b000, 12'hFFD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b000, 12'hFFE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b000, 12'hFFF} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h000} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h003} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'h004} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h005} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h007} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h008} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'h009} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h00B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h00C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h00D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h00E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h00F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h011} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h013} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h014} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h015} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h017} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b001, 12'h018} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h019} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h01B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h01D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h01F} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'h021} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h022} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h023} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h024} : s_CHIP_26B_45133_reg = 8'h48;
         {3'b001, 12'h025} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h027} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h028} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h029} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h02B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h02D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h02E} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b001, 12'h02F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h031} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h032} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h033} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b001, 12'h034} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'h035} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h037} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h039} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h03A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h03B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h03C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b001, 12'h03D} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'h03F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h041} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h042} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h043} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h045} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h047} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h049} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h04A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h04B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h04D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h04E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h04F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h051} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h053} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h055} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h056} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h057} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h058} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h059} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h05B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h05D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h05F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h060} : s_CHIP_26B_45133_reg = 8'h97;
         {3'b001, 12'h061} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h062} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h063} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h064} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b001, 12'h065} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h067} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h068} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h069} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h06B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h06C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h06D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h06F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h070} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b001, 12'h071} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h073} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h075} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h077} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h078} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h079} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h07B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h07C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h07D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h07F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h080} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h081} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h083} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h084} : s_CHIP_26B_45133_reg = 8'hE4;
         {3'b001, 12'h085} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h087} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h088} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h089} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h08B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h08D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h08F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h090} : s_CHIP_26B_45133_reg = 8'h3F;
         {3'b001, 12'h091} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h092} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h093} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h094} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h095} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h096} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h097} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b001, 12'h098} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h099} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'h09A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h09B} : s_CHIP_26B_45133_reg = 8'h42;
         {3'b001, 12'h09C} : s_CHIP_26B_45133_reg = 8'hA7;
         {3'b001, 12'h09D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h09F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h0A0} : s_CHIP_26B_45133_reg = 8'hA7;
         {3'b001, 12'h0A1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h0A3} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h0A4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h0A5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h0A6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h0A7} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h0A8} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h0AA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h0AB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h0AC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h0AD} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h0AF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h0B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h0B3} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h0B5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h0B7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'h0B9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h0BA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h0BB} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b001, 12'h0BC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h0BD} : s_CHIP_26B_45133_reg = 8'hB4;
         {3'b001, 12'h0BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h0C0} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h0C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h0C3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h0C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h0C7} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h0C9} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b001, 12'h0CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h0CD} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'h0CE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h0CF} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h0D1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h0D2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h0D3} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b001, 12'h0D4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h0D5} : s_CHIP_26B_45133_reg = 8'hB4;
         {3'b001, 12'h0D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h0D8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h0D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h0DB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h0DD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h0DE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h0DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h0E0} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h0E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h0E3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h0E4} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h0E5} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h0E7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h0E9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'h0EA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h0EB} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'h0EC} : s_CHIP_26B_45133_reg = 8'h38;
         {3'b001, 12'h0ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h0EE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h0EF} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h0F1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h0F3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h0F4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h0F5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h0F7} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'h0F8} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b001, 12'h0F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h0FA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h0FB} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h0FC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h0FD} : s_CHIP_26B_45133_reg = 8'hB4;
         {3'b001, 12'h0FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h100} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h101} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h103} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h104} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b001, 12'h105} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h107} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h109} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h10A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h10B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h10D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h10F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h110} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h111} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h112} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h113} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b001, 12'h114} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h115} : s_CHIP_26B_45133_reg = 8'hB4;
         {3'b001, 12'h117} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h118} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h119} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h11B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h11C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h11D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h11E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h11F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h121} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h122} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h123} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h124} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b001, 12'h125} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h126} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h127} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h128} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h129} : s_CHIP_26B_45133_reg = 8'hB4;
         {3'b001, 12'h12B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h12C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h12D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h12E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h12F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b001, 12'h131} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h133} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h134} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h135} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h137} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h139} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h13B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h13D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h13E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h13F} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h140} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h141} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h142} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h143} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h144} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h145} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h146} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'h147} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b001, 12'h149} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h14B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h14D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h14E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h14F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h151} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h153} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h154} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b001, 12'h155} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h157} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h158} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b001, 12'h159} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h15B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h15C} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h15D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h15F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h161} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h163} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h165} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h167} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h168} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b001, 12'h169} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h16A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h16B} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b001, 12'h16C} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b001, 12'h16D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h16F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h170} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h171} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h173} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h174} : s_CHIP_26B_45133_reg = 8'hC4;
         {3'b001, 12'h175} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h177} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h178} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h179} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h17B} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b001, 12'h17C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h17D} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h17F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h180} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b001, 12'h181} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h183} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h184} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h185} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h187} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h188} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h189} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h18B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h18C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h18D} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h18F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h190} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h191} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h193} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h194} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h195} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h197} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h198} : s_CHIP_26B_45133_reg = 8'hFC;
         {3'b001, 12'h199} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h19A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h19B} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b001, 12'h19D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h19F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h1A0} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b001, 12'h1A1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h1A3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h1A4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h1A5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h1A7} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h1A8} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b001, 12'h1AB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h1AC} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b001, 12'h1AD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h1AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h1B0} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b001, 12'h1B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1B3} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'h1B4} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b001, 12'h1B5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1B7} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'h1B8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h1B9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h1BB} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'h1BD} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h1BF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h1C0} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h1C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1C3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h1C4} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h1C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1C7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h1C8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h1C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1CB} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h1CC} : s_CHIP_26B_45133_reg = 8'h1F;
         {3'b001, 12'h1CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1CF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h1D0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h1D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1D3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h1D4} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h1D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1D7} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h1D8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h1D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1DB} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h1DC} : s_CHIP_26B_45133_reg = 8'hC2;
         {3'b001, 12'h1DD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h1DF} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h1E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1E2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h1E3} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h1E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1E7} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h1EA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h1EB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h1EC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h1ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1EF} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h1F0} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h1F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1F3} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h1F4} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h1F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1F7} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h1F8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h1F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1FB} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h1FC} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h1FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h1FF} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h200} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h201} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h203} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h204} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h205} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h207} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h208} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b001, 12'h209} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h20B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h20C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h20D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h20F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h210} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h211} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h213} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h214} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h215} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h216} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h217} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h218} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h219} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h21B} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b001, 12'h21C} : s_CHIP_26B_45133_reg = 8'hC7;
         {3'b001, 12'h21D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h21F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h221} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h222} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h223} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h225} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h227} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h229} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h22B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h22C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h22D} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'h22E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h22F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h230} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h231} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h233} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b001, 12'h234} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h235} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h237} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b001, 12'h238} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b001, 12'h239} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h23B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b001, 12'h23C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'h23D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h23F} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b001, 12'h241} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h243} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h244} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h245} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h247} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b001, 12'h248} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h249} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h24B} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b001, 12'h24C} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h24D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h24E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h24F} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b001, 12'h250} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'h251} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h253} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b001, 12'h254} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b001, 12'h255} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h257} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h258} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'h259} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h25A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h25B} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b001, 12'h25C} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b001, 12'h25D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h25F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h260} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h261} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h263} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b001, 12'h264} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h265} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h266} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h267} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'h268} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b001, 12'h269} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h26A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h26B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h26C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h26D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h26F} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h270} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h271} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h273} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h274} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h277} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h279} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h27A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h27B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h27C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h27D} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b001, 12'h27F} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b001, 12'h280} : s_CHIP_26B_45133_reg = 8'hC4;
         {3'b001, 12'h281} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h283} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h285} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h286} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h287} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h288} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h289} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h28B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h28D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h28F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h290} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h291} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'h292} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h293} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h295} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h297} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h298} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h299} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h29B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h29C} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b001, 12'h29E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h29F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h2A0} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h2A1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h2A3} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h2A4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2A8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2A9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h2AB} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h2AD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h2B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h2B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2B4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2B5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2B8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h2BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2BC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h2BD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h2BF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h2C0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2C1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2C4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2C8} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2C9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h2CB} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'h2CC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h2CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h2CF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h2D0} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h2D1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h2D2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h2D3} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b001, 12'h2D4} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h2D5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h2D6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h2D7} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b001, 12'h2D8} : s_CHIP_26B_45133_reg = 8'hA4;
         {3'b001, 12'h2D9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2DA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h2DB} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b001, 12'h2DC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2DD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2E0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2E4} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h2E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h2E7} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b001, 12'h2E8} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2E9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h2EB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h2EC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2ED} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h2EF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h2F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h2F3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h2F4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h2F5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h2F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h2F9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h2FB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'h2FC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'h2FD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h2FE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h2FF} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h300} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h301} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h303} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h304} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h305} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h307} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h309} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h30B} : s_CHIP_26B_45133_reg = 8'h38;
         {3'b001, 12'h30C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h30D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h30F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h310} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h311} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h313} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h314} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h315} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h317} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h318} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h319} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h31B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h31C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h31F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h320} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h321} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h323} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b001, 12'h324} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h325} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h326} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h327} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'h328} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h329} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h32B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h32C} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h32D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h32F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h330} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h333} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h334} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h335} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h337} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h338} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'h33A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h33B} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b001, 12'h33C} : s_CHIP_26B_45133_reg = 8'hD4;
         {3'b001, 12'h33F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h340} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h341} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h343} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h344} : s_CHIP_26B_45133_reg = 8'hD4;
         {3'b001, 12'h345} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h347} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h348} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h349} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h34B} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'h34D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h34F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h350} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h351} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h352} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h353} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b001, 12'h354} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h355} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b001, 12'h356} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h357} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b001, 12'h358} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h359} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h35B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h35C} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h35D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h35F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h361} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h363} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h364} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h365} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h366} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h367} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h369} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h36B} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b001, 12'h36D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h36E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h36F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h370} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b001, 12'h371} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h373} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'h375} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h376} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h377} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h378} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h379} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h37B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h37E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h37F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h381} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h382} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h383} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h384} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h385} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h387} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h388} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h389} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h38A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h38B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h38C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h38D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h38F} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b001, 12'h390} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b001, 12'h391} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h393} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b001, 12'h394} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h396} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h397} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h399} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h39B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h39C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h39D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h39F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h3A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h3A2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h3A3} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b001, 12'h3A4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h3A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3A6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h3A7} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b001, 12'h3A8} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h3A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3AB} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h3AC} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h3AD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h3AF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h3B0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3B1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h3B5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h3B7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h3B8} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b001, 12'h3B9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3BB} : s_CHIP_26B_45133_reg = 8'h25;
         {3'b001, 12'h3BC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h3BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h3BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3BF} : s_CHIP_26B_45133_reg = 8'hFB;
         {3'b001, 12'h3C0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h3C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h3C2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3C3} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b001, 12'h3C4} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h3C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h3C6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3C7} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b001, 12'h3C8} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h3C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h3CB} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'h3CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h3CF} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b001, 12'h3D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h3D3} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h3D4} : s_CHIP_26B_45133_reg = 8'hE4;
         {3'b001, 12'h3D7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h3D8} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h3DB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h3DC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h3DD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h3DF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h3E0} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b001, 12'h3E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3E3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h3E5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h3E6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h3E7} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h3E8} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3EA} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h3EB} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h3EC} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b001, 12'h3ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h3EF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h3F0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h3F1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h3F3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h3F4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h3F5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h3F7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h3F8} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b001, 12'h3F9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h3FB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h3FC} : s_CHIP_26B_45133_reg = 8'hF5;
         {3'b001, 12'h3FE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h3FF} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h400} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h401} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h402} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h403} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h404} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h405} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h407} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h408} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h409} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h40B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h40C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h40D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h40F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h410} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h411} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h412} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h413} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b001, 12'h414} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b001, 12'h415} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h417} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h418} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h419} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h41A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h41B} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h41C} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b001, 12'h41F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h420} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h421} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h422} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h423} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b001, 12'h425} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h427} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h428} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h429} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h42B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h42C} : s_CHIP_26B_45133_reg = 8'hF5;
         {3'b001, 12'h42E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h42F} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h430} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h431} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h432} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h433} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b001, 12'h434} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h436} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h437} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h438} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h439} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h43B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h43C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h43D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h43F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h440} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h441} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h443} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h444} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b001, 12'h447} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h448} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b001, 12'h449} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h44B} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b001, 12'h44C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h44D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h44F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h450} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b001, 12'h451} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h453} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b001, 12'h455} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h456} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h457} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h458} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h459} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h45B} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b001, 12'h45C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h45D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h45F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h461} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h462} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h463} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b001, 12'h464} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'h465} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h467} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h468} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h469} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h46B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h46C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b001, 12'h46D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h46E} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b001, 12'h46F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h471} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h472} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h473} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h475} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h477} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b001, 12'h479} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h47A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h47B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h47D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h47F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'h480} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h481} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h482} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h483} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h485} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h486} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h487} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h488} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h48B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h48D} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b001, 12'h48F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h491} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h492} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h493} : s_CHIP_26B_45133_reg = 8'h67;
         {3'b001, 12'h494} : s_CHIP_26B_45133_reg = 8'h95;
         {3'b001, 12'h495} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h496} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h497} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b001, 12'h498} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h499} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h49B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h49D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h49E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h49F} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h4A0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4A3} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h4A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h4A6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h4A7} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h4A8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h4AC} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'h4AD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h4AE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h4AF} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h4B0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4B1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4B2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h4B3} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h4B4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4B5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4B6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h4B7} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h4B8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h4B9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4BA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h4BB} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h4BC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4BD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4BE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h4BF} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h4C0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4C1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4C2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h4C3} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h4C4} : s_CHIP_26B_45133_reg = 8'h75;
         {3'b001, 12'h4C5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4C6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h4C7} : s_CHIP_26B_45133_reg = 8'h67;
         {3'b001, 12'h4C8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4C9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h4CB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'h4CD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h4CE} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h4CF} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h4D0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4D1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4D3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h4D4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4D5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4D6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h4D7} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h4D8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4D9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4DA} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h4DB} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h4DC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4DD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4DE} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h4DF} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h4E0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4E2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h4E3} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h4E4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4E6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h4E7} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h4E8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h4E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h4ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h4EF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h4F0} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h4F3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h4F5} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b001, 12'h4F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h4F8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h4F9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h4FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h4FC} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h4FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h4FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h500} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h501} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h503} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h507} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h508} : s_CHIP_26B_45133_reg = 8'hF8;
         {3'b001, 12'h509} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h50B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h50C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h50D} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h50E} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b001, 12'h50F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h510} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h511} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h513} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h515} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h516} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b001, 12'h517} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h518} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h519} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h51A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h51B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h51C} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b001, 12'h51D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h51F} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b001, 12'h521} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h523} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h525} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h526} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h527} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h528} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h529} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h52B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h52D} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h52E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h52F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h531} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h533} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h535} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h536} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h537} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'h538} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h539} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h53A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h53B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h53C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h53D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h53E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h53F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'h540} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h541} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h543} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b001, 12'h544} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h545} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h547} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h549} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h54A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h54B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h54D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h54F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h550} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h551} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h553} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h554} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h555} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h557} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b001, 12'h558} : s_CHIP_26B_45133_reg = 8'hF5;
         {3'b001, 12'h55B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h55D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h55E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h55F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h560} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h561} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h563} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h565} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h567} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h568} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h56B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h56D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h56E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h56F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h571} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h573} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h574} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h575} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h577} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h578} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b001, 12'h579} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'h57B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b001, 12'h57C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h57F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h580} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h581} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h583} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h584} : s_CHIP_26B_45133_reg = 8'hC5;
         {3'b001, 12'h587} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h588} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h589} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h58A} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b001, 12'h58B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h58C} : s_CHIP_26B_45133_reg = 8'h25;
         {3'b001, 12'h58E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h58F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h591} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h592} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h593} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h595} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h596} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b001, 12'h597} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h598} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h59A} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b001, 12'h59B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h59C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h59D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h59E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h59F} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b001, 12'h5A0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h5A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5A3} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'h5A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5A7} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b001, 12'h5A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5AB} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h5AC} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h5AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5AF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h5B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5B3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h5B4} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h5B5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h5B7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h5B8} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h5B9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h5BB} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h5BC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h5BD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h5BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h5C1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h5C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h5C4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h5C5} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h5C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h5C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5CA} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b001, 12'h5CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h5CC} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h5CD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h5CE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h5CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h5D0} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h5D2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h5D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h5D4} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h5D5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h5D7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h5D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5DA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h5DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h5DC} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h5DD} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h5DF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h5E0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h5E1} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'h5E3} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'h5E4} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h5E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5E7} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h5E8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h5E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5EB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h5EC} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h5ED} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h5EF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h5F0} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b001, 12'h5F1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h5F3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h5F4} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h5F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5F7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h5F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5FB} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'h5FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h5FF} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'h601} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h603} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'h604} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h605} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h607} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'h608} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h609} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h60B} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h60C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h60D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h60F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h610} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h611} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h613} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h614} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h615} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h617} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h618} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h619} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h61B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h61F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h620} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h621} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h623} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h624} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b001, 12'h625} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h627} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'h628} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h62B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h62C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h62D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h62F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h630} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h631} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h633} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h634} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h635} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h637} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h638} : s_CHIP_26B_45133_reg = 8'hE4;
         {3'b001, 12'h639} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h63B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h63C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h63F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h640} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h643} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h644} : s_CHIP_26B_45133_reg = 8'hC5;
         {3'b001, 12'h645} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h647} : s_CHIP_26B_45133_reg = 8'hFB;
         {3'b001, 12'h649} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h64B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h64C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h64D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h64F} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'h650} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h651} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h653} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'h654} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h657} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h658} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h659} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h65B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h65C} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h65D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h65F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h660} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h661} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h663} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h664} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h665} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h667} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h668} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h66B} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'h66C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h66D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h66F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h670} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h671} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h673} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h675} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h677} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h679} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h67B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h67D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h67F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h680} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h681} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h683} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h684} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h685} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h687} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h688} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h689} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h68B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h68C} : s_CHIP_26B_45133_reg = 8'hA5;
         {3'b001, 12'h68D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h68F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h690} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'h691} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h693} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h694} : s_CHIP_26B_45133_reg = 8'h15;
         {3'b001, 12'h695} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h697} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b001, 12'h698} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h699} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h69A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h69B} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h69C} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b001, 12'h69D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h69E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h69F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h6A0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h6A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h6A2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h6A3} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h6A5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h6A6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h6A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h6A8} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h6A9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h6AB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h6AC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h6AD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h6AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h6B0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h6B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h6B3} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b001, 12'h6B4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h6B5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h6B7} : s_CHIP_26B_45133_reg = 8'h3D;
         {3'b001, 12'h6B8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h6B9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h6BB} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b001, 12'h6BC} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'h6BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h6BF} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'h6C0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h6C1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h6C3} : s_CHIP_26B_45133_reg = 8'h3D;
         {3'b001, 12'h6C4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h6C5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h6C7} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b001, 12'h6C8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h6C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h6CB} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b001, 12'h6CC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h6CD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h6CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h6D0} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h6D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h6D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h6D7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h6D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h6DB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'h6DC} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h6DD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h6DF} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b001, 12'h6E0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h6E3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'h6E4} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h6E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h6E7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h6E8} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h6E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h6EB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h6EC} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b001, 12'h6EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h6F0} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h6F1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h6F3} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h6F4} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h6F5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h6F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h6F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h6FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h6FE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h6FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h700} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h701} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h703} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h704} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h705} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h707} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h708} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h709} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h70B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h70D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h70F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h711} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h713} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h715} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h716} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h717} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h718} : s_CHIP_26B_45133_reg = 8'hC5;
         {3'b001, 12'h71B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h71D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h71F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h720} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h721} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h723} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h727} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h728} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h729} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h72B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h72C} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h72D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h72F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h730} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h731} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h733} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h734} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h735} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h736} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h737} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h738} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h73B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h73C} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h73D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h73F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h740} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h743} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h744} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h745} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h747} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h748} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h749} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h74B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h74C} : s_CHIP_26B_45133_reg = 8'hC6;
         {3'b001, 12'h74D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h74F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h751} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h752} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h753} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h754} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h755} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h756} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h757} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h758} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h759} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h75A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h75B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h75C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h75D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h75F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h760} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h761} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h763} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h765} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h767} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h768} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h769} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h76B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h76C} : s_CHIP_26B_45133_reg = 8'hB6;
         {3'b001, 12'h76F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h771} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h772} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h773} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h774} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h775} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h776} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h777} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h778} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h779} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h77B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h77C} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h77D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h77F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h781} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h783} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b001, 12'h785} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h787} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b001, 12'h788} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h789} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h78B} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'h78C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h78D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h78F} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h790} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h791} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h793} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'h794} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h795} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h797} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h798} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h79A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h79B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h79C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h79D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h79F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h7A2} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b001, 12'h7A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7A4} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h7A5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h7A6} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h7A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7A8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h7AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h7AE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h7AF} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h7B0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h7B1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h7B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7B4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h7B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h7BA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h7BB} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h7BC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h7BD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h7BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7C0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h7C2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'h7C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7C4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h7C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h7C6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h7C7} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h7C8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h7C9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h7CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7CC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h7CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7D0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h7D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h7D3} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h7D4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h7D5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h7D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7D8} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h7D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h7DB} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h7DC} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h7DD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h7DF} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h7E0} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h7E1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h7E3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h7E4} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h7E5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h7E6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h7E7} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h7E8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h7E9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h7EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7EC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h7EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h7F2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h7F3} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b001, 12'h7F4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h7F5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h7F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h7F8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h7F9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h7FB} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h7FC} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h7FD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h7FF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h800} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h801} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h802} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h803} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h804} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h805} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h807} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h808} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h809} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h80B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h80C} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h80D} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b001, 12'h80E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h80F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h810} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h813} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h814} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h815} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h816} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h817} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h818} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h819} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h81A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h81B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h81C} : s_CHIP_26B_45133_reg = 8'hD6;
         {3'b001, 12'h81D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h81F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h820} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h821} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h823} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'h824} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h827} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h828} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h829} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h82B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h82C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h82F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h831} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h833} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b001, 12'h835} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h836} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h837} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h838} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h839} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h83B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h83C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h83D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h83F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h840} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h841} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h843} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h844} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h845} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h847} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b001, 12'h849} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h84A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h84B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h84C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h84D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h84F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h850} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h851} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h853} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h854} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h857} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h858} : s_CHIP_26B_45133_reg = 8'h56;
         {3'b001, 12'h859} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h85B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h85C} : s_CHIP_26B_45133_reg = 8'hF5;
         {3'b001, 12'h85F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h860} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h861} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h862} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h863} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h865} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h867} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h868} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h869} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h86B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h86C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h86F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'h870} : s_CHIP_26B_45133_reg = 8'h56;
         {3'b001, 12'h871} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h872} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h873} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h874} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h875} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h876} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h877} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h878} : s_CHIP_26B_45133_reg = 8'hB6;
         {3'b001, 12'h87B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h87C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h87D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h87F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h880} : s_CHIP_26B_45133_reg = 8'hD6;
         {3'b001, 12'h881} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h882} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h883} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b001, 12'h884} : s_CHIP_26B_45133_reg = 8'hC6;
         {3'b001, 12'h887} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h889} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h88A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h88B} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b001, 12'h88C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h88D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h88F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h890} : s_CHIP_26B_45133_reg = 8'hD6;
         {3'b001, 12'h891} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h892} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h893} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b001, 12'h894} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h895} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h896} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h897} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b001, 12'h899} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h89B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h89C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h89D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h89F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h8A0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h8A3} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h8A4} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h8A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h8A7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h8A8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h8A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h8AB} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'h8AC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h8AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h8AF} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'h8B0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h8B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h8B3} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'h8B4} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h8B5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h8B7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h8B8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h8B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h8BB} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'h8BC} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h8BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h8BF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h8C1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h8C2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h8C3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h8C4} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'h8C5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h8C7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h8C8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8C9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8CA} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h8CB} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h8CC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8CD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8CE} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h8CF} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h8D0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8D1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8D2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h8D3} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h8D4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8D5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8D6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h8D7} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h8D8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8D9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8DA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h8DB} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h8DC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8DD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8DE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h8DF} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h8E0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8E2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h8E3} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h8E4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8E6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h8E7} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h8E8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8EA} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h8EB} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h8EC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8EE} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h8EF} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h8F0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8F1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8F2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h8F3} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h8F4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8F5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8F6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h8F7} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h8F8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h8F9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8FA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h8FB} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h8FC} : s_CHIP_26B_45133_reg = 8'hA6;
         {3'b001, 12'h8FD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h8FE} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h8FF} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'h900} : s_CHIP_26B_45133_reg = 8'h56;
         {3'b001, 12'h901} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h902} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h903} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h904} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h907} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h908} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h90A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h90B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h90C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h90E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h90F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h910} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h912} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h913} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h914} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h916} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h917} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h918} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h91A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h91B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h91C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h91E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h91F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h920} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h922} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h923} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h924} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h926} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h927} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h928} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h929} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h92B} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'h92C} : s_CHIP_26B_45133_reg = 8'hD6;
         {3'b001, 12'h92F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h930} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h933} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h934} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h935} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h937} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h938} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b001, 12'h93A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'h93B} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b001, 12'h93D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h93F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'h940} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h941} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h943} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h944} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h945} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h947} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h948} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h949} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h94B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h94C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'h94D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h94F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h950} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h951} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h953} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h954} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'h955} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h957} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b001, 12'h958} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h959} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h95B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h95C} : s_CHIP_26B_45133_reg = 8'hD6;
         {3'b001, 12'h95F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h960} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h961} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h963} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h964} : s_CHIP_26B_45133_reg = 8'hD5;
         {3'b001, 12'h965} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h967} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h968} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h969} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h96B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'h96C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h96D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h96F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h970} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'h973} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h974} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h975} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h977} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h978} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'h979} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h97A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h97B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h97D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h97F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'h980} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'h981} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h983} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h984} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h985} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h987} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'h988} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b001, 12'h989} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h98B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b001, 12'h98C} : s_CHIP_26B_45133_reg = 8'hC5;
         {3'b001, 12'h98F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'h990} : s_CHIP_26B_45133_reg = 8'hE6;
         {3'b001, 12'h992} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'h993} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h995} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h997} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h998} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b001, 12'h99B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h99D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h99E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h99F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h9A0} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'h9A1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h9A3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'h9A4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h9A5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'h9A7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'h9A8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h9A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h9AB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'h9AD} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'h9AE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h9AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h9B0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h9B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h9B3} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b001, 12'h9B4} : s_CHIP_26B_45133_reg = 8'hD6;
         {3'b001, 12'h9B5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h9B7} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'h9B8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h9B9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h9BB} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h9BC} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b001, 12'h9BD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h9BF} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b001, 12'h9C0} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b001, 12'h9C1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h9C3} : s_CHIP_26B_45133_reg = 8'hEE;
         {3'b001, 12'h9C4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h9C5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'h9C7} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'h9C8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'h9C9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h9CB} : s_CHIP_26B_45133_reg = 8'hEE;
         {3'b001, 12'h9CC} : s_CHIP_26B_45133_reg = 8'hFC;
         {3'b001, 12'h9CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h9CF} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b001, 12'h9D0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'h9D1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h9D3} : s_CHIP_26B_45133_reg = 8'hFB;
         {3'b001, 12'h9D4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'h9D5} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b001, 12'h9D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h9D9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'h9DB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'h9DC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h9E0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h9E4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'h9E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h9EA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'h9EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h9ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h9EF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h9F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h9F2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'h9F3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'h9F4} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h9F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'h9F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'h9F8} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'h9F9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'h9FB} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b001, 12'h9FC} : s_CHIP_26B_45133_reg = 8'h56;
         {3'b001, 12'h9FD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'h9FF} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hA00} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hA01} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hA03} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hA04} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hA05} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b001, 12'hA06} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hA07} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b001, 12'hA09} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hA0B} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b001, 12'hA0C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hA0D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hA0E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hA0F} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b001, 12'hA10} : s_CHIP_26B_45133_reg = 8'hB7;
         {3'b001, 12'hA11} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hA13} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b001, 12'hA14} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hA15} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hA17} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hA18} : s_CHIP_26B_45133_reg = 8'hB6;
         {3'b001, 12'hA19} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hA1A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hA1B} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b001, 12'hA1C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hA1D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hA1F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hA20} : s_CHIP_26B_45133_reg = 8'hB6;
         {3'b001, 12'hA21} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hA23} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b001, 12'hA25} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA27} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'hA28} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hA29} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA2B} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'hA2C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hA2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA2F} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'hA30} : s_CHIP_26B_45133_reg = 8'h56;
         {3'b001, 12'hA33} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hA34} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hA37} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hA39} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA3B} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'hA3C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hA3D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA3F} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hA40} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hA41} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA43} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'hA44} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hA45} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA47} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hA48} : s_CHIP_26B_45133_reg = 8'hA6;
         {3'b001, 12'hA4B} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'hA4D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA4F} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'hA50} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hA51} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA53} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'hA54} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hA55} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA57} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'hA58} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hA59} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA5B} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hA5D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA5F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hA60} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hA61} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA63} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b001, 12'hA64} : s_CHIP_26B_45133_reg = 8'hB6;
         {3'b001, 12'hA67} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b001, 12'hA69} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA6B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hA6C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hA6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA6F} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b001, 12'hA70} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hA71} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b001, 12'hA73} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b001, 12'hA75} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hA76} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hA77} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b001, 12'hA79} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA7A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hA7B} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'hA7C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hA7D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hA7F} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b001, 12'hA80} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hA81} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hA83} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hA84} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hA85} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA88} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hA89} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hA8A} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA8B} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'hA8C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hA8D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA8F} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hA90} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b001, 12'hA91} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hA93} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'hA94} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hA95} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA97} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b001, 12'hA99} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA9A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hA9B} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b001, 12'hA9D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hA9F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'hAA0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hAA1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAA3} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b001, 12'hAA4} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hAA5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAA7} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hAA8} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hAA9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hAAB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hAAC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hAAF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hAB0} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hAB1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAB3} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hAB4} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hAB7} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hAB8} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hAB9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hABB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hABC} : s_CHIP_26B_45133_reg = 8'h97;
         {3'b001, 12'hABF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hAC0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hAC1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAC3} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b001, 12'hAC4} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hAC5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hAC6} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAC7} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hAC8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hAC9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hACB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hACD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hACE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hACF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b001, 12'hAD0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hAD2} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAD3} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b001, 12'hAD4} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAD5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAD7} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b001, 12'hAD8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hAD9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hADB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hADD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hADF} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b001, 12'hAE1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAE3} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b001, 12'hAE4} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'hAE5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hAE7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hAE8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hAE9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hAEB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hAEC} : s_CHIP_26B_45133_reg = 8'hE6;
         {3'b001, 12'hAED} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hAEF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hAF1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hAF3} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hAF4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hAF7} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hAF8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hAF9} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b001, 12'hAFB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hAFD} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hAFE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hAFF} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b001, 12'hB01} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB02} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hB03} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b001, 12'hB05} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB06} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hB07} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b001, 12'hB08} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hB09} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hB0A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'hB0B} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hB0D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB0E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hB0F} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b001, 12'hB11} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hB13} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'hB15} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hB16} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hB17} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'hB19} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB1B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hB1D} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hB1F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'hB20} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'hB21} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hB22} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hB23} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b001, 12'hB24} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hB25} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB27} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hB28} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hB29} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hB2A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hB2B} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hB2C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hB2F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hB30} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hB31} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB33} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'hB34} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hB35} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hB37} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'hB38} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hB39} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b001, 12'hB3B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hB3D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hB3E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hB3F} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'hB41} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB43} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'hB44} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hB45} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hB46} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b001, 12'hB47} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hB49} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB4B} : s_CHIP_26B_45133_reg = 8'h67;
         {3'b001, 12'hB4D} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hB4F} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'hB51} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hB52} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hB53} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b001, 12'hB54} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hB56} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hB57} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hB58} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hB59} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB5B} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hB5C} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hB5F} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hB61} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB62} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hB63} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hB65} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB67} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hB69} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB6B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hB6C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hB6D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hB6F} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b001, 12'hB70} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hB71} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hB73} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hB74} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hB75} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB77} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hB78} : s_CHIP_26B_45133_reg = 8'hB6;
         {3'b001, 12'hB79} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hB7C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB7D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB7F} : s_CHIP_26B_45133_reg = 8'h77;
         {3'b001, 12'hB80} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hB81} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hB83} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b001, 12'hB84} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b001, 12'hB85} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hB87} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hB88} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hB89} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB8B} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hB8C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hB8D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB8F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hB90} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hB91} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hB93} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hB94} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hB95} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hB97} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hB98} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hB99} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB9B} : s_CHIP_26B_45133_reg = 8'h1C;
         {3'b001, 12'hB9C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hB9D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hB9F} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hBA0} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hBA1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hBA3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hBA4} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hBA5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBA7} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b001, 12'hBA8} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hBA9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBAB} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'hBAC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hBAD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBAF} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'hBB0} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'hBB1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBB3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hBB4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hBB5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBB7} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hBB8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hBB9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBBB} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hBBD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hBBF} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b001, 12'hBC1} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hBC3} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hBC4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hBC5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBC6} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hBC8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hBC9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hBCA} : s_CHIP_26B_45133_reg = 8'h98;
         {3'b001, 12'hBCB} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBCC} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hBCD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBCF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hBD1} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hBD2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hBD3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hBD4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hBD5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBD6} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hBD8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hBD9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hBDA} : s_CHIP_26B_45133_reg = 8'h98;
         {3'b001, 12'hBDB} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBDC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hBDD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBDE} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hBE0} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hBE1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hBE2} : s_CHIP_26B_45133_reg = 8'h98;
         {3'b001, 12'hBE3} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'hBE4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'hBE5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBE7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hBE8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hBE9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBEB} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hBEC} : s_CHIP_26B_45133_reg = 8'hB7;
         {3'b001, 12'hBED} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hBEF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hBF0} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hBF1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hBF3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hBF4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hBF5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hBF7} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'hBF8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hBF9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hBFB} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b001, 12'hBFC} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hBFD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hBFE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hBFF} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hC00} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hC03} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hC04} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hC05} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC07} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b001, 12'hC09} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC0A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hC0B} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b001, 12'hC0D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC0F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'hC10} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hC13} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hC15} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC16} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hC17} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hC19} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC1B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hC1C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hC1D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC1F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hC21} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC23} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hC24} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hC25} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hC27} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b001, 12'hC28} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hC29} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hC2B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hC2C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hC2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC2F} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hC30} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hC31} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hC32} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hC33} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hC34} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hC35} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC37} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b001, 12'hC38} : s_CHIP_26B_45133_reg = 8'hF7;
         {3'b001, 12'hC39} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hC3B} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b001, 12'hC3C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'hC3D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC3F} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'hC40} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hC41} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC43} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hC44} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hC45} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hC47} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hC48} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hC49} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hC4B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hC4C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hC4D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hC4F} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hC50} : s_CHIP_26B_45133_reg = 8'h57;
         {3'b001, 12'hC51} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hC53} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b001, 12'hC54} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hC55} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hC57} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hC58} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hC59} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hC5B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hC5C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hC5D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hC5F} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hC60} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hC61} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hC63} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hC64} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hC67} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hC69} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC6B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hC6C} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hC6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC6F} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'hC70} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hC71} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC73} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'hC74} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hC75} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC77} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hC78} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hC79} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC7B} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hC7D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC7F} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'hC80} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'hC81} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hC83} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hC84} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hC85} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC86} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hC87} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hC88} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hC89} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hC8A} : s_CHIP_26B_45133_reg = 8'h88;
         {3'b001, 12'hC8B} : s_CHIP_26B_45133_reg = 8'hC4;
         {3'b001, 12'hC8C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hC8D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC8E} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hC8F} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hC90} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hC91} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hC92} : s_CHIP_26B_45133_reg = 8'hA8;
         {3'b001, 12'hC93} : s_CHIP_26B_45133_reg = 8'hC4;
         {3'b001, 12'hC95} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC97} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hC99} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hC9B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hC9C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hC9D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hC9E} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hC9F} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hCA0} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hCA1} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hCA2} : s_CHIP_26B_45133_reg = 8'hA8;
         {3'b001, 12'hCA3} : s_CHIP_26B_45133_reg = 8'hC4;
         {3'b001, 12'hCA4} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hCA5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hCA7} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hCA8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hCA9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hCAB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hCAD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCAE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hCAF} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b001, 12'hCB0} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'hCB1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCB3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'hCB4} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hCB5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCB7} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hCB8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hCB9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCBB} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hCBC} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hCBD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hCBF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hCC0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'hCC1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCC3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hCC4} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCC7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hCC8} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'hCC9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCCB} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'hCCC} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hCCD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCCF} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b001, 12'hCD0} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hCD3} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hCD5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCD7} : s_CHIP_26B_45133_reg = 8'h7E;
         {3'b001, 12'hCD8} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b001, 12'hCD9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCDB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hCDC} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hCDD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCDF} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b001, 12'hCE1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCE3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hCE4} : s_CHIP_26B_45133_reg = 8'h87;
         {3'b001, 12'hCE7} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hCE8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hCE9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hCEB} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b001, 12'hCEC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hCED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCEF} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hCF0} : s_CHIP_26B_45133_reg = 8'h56;
         {3'b001, 12'hCF1} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'hCF3} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b001, 12'hCF5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCF7} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b001, 12'hCF8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hCF9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hCFB} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'hCFC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hCFD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hCFF} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b001, 12'hD00} : s_CHIP_26B_45133_reg = 8'hB7;
         {3'b001, 12'hD01} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b001, 12'hD03} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b001, 12'hD04} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD05} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD07} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hD08} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hD09} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hD0B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hD0C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hD0D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hD0F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hD12} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hD13} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hD15} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD16} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hD17} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b001, 12'hD18} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hD19} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hD1B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hD1C} : s_CHIP_26B_45133_reg = 8'h97;
         {3'b001, 12'hD1D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hD1F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hD20} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hD21} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD23} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b001, 12'hD25} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD26} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hD27} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b001, 12'hD29} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b001, 12'hD2B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b001, 12'hD2D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hD2E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hD2F} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b001, 12'hD31} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD32} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hD33} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b001, 12'hD34} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hD35} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD36} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hD37} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b001, 12'hD38} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hD39} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD3A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hD3B} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b001, 12'hD3D} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b001, 12'hD3F} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'hD41} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hD43} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'hD45} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD47} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b001, 12'hD48} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b001, 12'hD4A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hD4B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hD4D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD4F} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b001, 12'hD51} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b001, 12'hD52} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hD53} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hD55} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hD57} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b001, 12'hD58} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b001, 12'hD59} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD5B} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b001, 12'hD5C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hD5D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD5F} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b001, 12'hD60} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hD61} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD65} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD67} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b001, 12'hD68} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hD69} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD6B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hD6C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b001, 12'hD6D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hD6F} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hD70} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hD71} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hD73} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hD74} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD75} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hD77} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b001, 12'hD78} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hD79} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hD7B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hD7C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b001, 12'hD7D} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b001, 12'hD7F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hD81} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b001, 12'hD82} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b001, 12'hD83} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b001, 12'hD85} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD87} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'hD88} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hD89} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hD8B} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b001, 12'hD8C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hD8D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hD8F} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b001, 12'hD91} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD92} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hD93} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b001, 12'hD94} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b001, 12'hD95} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hD97} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hD9A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hD9B} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hD9C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hD9F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hDA0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hDA4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hDA8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hDAC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hDB0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hDB4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hDB8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hDBC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hDC1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDC3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDC4} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hDC5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDC7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDC8} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b001, 12'hDC9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDCB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDCC} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b001, 12'hDCD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDCF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDD0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hDD1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDD3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDD4} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hDD5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDD7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDD8} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b001, 12'hDD9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDDB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDDD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDDF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDE0} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hDE1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDE3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDE4} : s_CHIP_26B_45133_reg = 8'h83;
         {3'b001, 12'hDE5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDE7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDE8} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b001, 12'hDE9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDEB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDEC} : s_CHIP_26B_45133_reg = 8'hA3;
         {3'b001, 12'hDED} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDEF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDF0} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hDF1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDF3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDF4} : s_CHIP_26B_45133_reg = 8'h83;
         {3'b001, 12'hDF5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDF7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDF8} : s_CHIP_26B_45133_reg = 8'hA3;
         {3'b001, 12'hDF9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDFB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hDFC} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hDFD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hDFF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hE00} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hE01} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE02} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE03} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE04} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hE05} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE06} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE07} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE08} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hE09} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE0A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE0C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hE0D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE0E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE0F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE10} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hE11} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE12} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE13} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hE15} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE16} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE17} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'hE18} : s_CHIP_26B_45133_reg = 8'h53;
         {3'b001, 12'hE19} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE1A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE1B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hE1C} : s_CHIP_26B_45133_reg = 8'h53;
         {3'b001, 12'hE1D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE1E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE1F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hE20} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hE21} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE22} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE23} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE24} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hE25} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE26} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE27} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE28} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hE29} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE2A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE2B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE2C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b001, 12'hE2D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE2E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE2F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE30} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hE31} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE32} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE33} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hE35} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE36} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE37} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b001, 12'hE38} : s_CHIP_26B_45133_reg = 8'h53;
         {3'b001, 12'hE39} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE3A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE3B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hE3C} : s_CHIP_26B_45133_reg = 8'h53;
         {3'b001, 12'hE3D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE3E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b001, 12'hE3F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hE40} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'hE43} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE44} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b001, 12'hE47} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hE48} : s_CHIP_26B_45133_reg = 8'h35;
         {3'b001, 12'hE4B} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b001, 12'hE4C} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b001, 12'hE4F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b001, 12'hE50} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hE51} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hE53} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hE54} : s_CHIP_26B_45133_reg = 8'hC7;
         {3'b001, 12'hE55} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE57} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b001, 12'hE58} : s_CHIP_26B_45133_reg = 8'hC5;
         {3'b001, 12'hE5B} : s_CHIP_26B_45133_reg = 8'h25;
         {3'b001, 12'hE5C} : s_CHIP_26B_45133_reg = 8'hC5;
         {3'b001, 12'hE5D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hE5F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hE60} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE61} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b001, 12'hE62} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hE63} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b001, 12'hE64} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'hE65} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b001, 12'hE66} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hE67} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b001, 12'hE68} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b001, 12'hE6B} : s_CHIP_26B_45133_reg = 8'h25;
         {3'b001, 12'hE6C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b001, 12'hE6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hE6F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hE70} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b001, 12'hE71} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b001, 12'hE73} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hE74} : s_CHIP_26B_45133_reg = 8'hC5;
         {3'b001, 12'hE77} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE78} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hE7C} : s_CHIP_26B_45133_reg = 8'hC5;
         {3'b001, 12'hE7F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hE80} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'hE83} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE84} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b001, 12'hE87} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b001, 12'hE88} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b001, 12'hE8B} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'hE8C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'hE8F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hE90} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b001, 12'hE93} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b001, 12'hE94} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hE97} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b001, 12'hE98} : s_CHIP_26B_45133_reg = 8'hD1;
         {3'b001, 12'hE9B} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'hE9C} : s_CHIP_26B_45133_reg = 8'hD1;
         {3'b001, 12'hE9F} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b001, 12'hEA0} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b001, 12'hEA3} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'hEA4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'hEA7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hEA8} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b001, 12'hEAB} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'hEAC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'hEAF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hEB0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b001, 12'hEB3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hEB4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hEB7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hEB8} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b001, 12'hEBB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hEBC} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b001, 12'hEBF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hEC1} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hEC2} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hEC3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hEC5} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hEC7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hEC8} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b001, 12'hECB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hECC} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b001, 12'hECF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hED0} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b001, 12'hED3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hED4} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b001, 12'hED6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hED7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hED8} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hEDA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hEDB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hEDC} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b001, 12'hEDF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hEE1} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hEE2} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hEE3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hEE5} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hEE7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hEE8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hEEA} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hEEB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hEEC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hEEE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hEEF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hEF0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hEF3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hEF4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hEF6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hEF7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b001, 12'hEF9} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hEFB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hEFC} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b001, 12'hEFF} : s_CHIP_26B_45133_reg = 8'h1F;
         {3'b001, 12'hF00} : s_CHIP_26B_45133_reg = 8'h52;
         {3'b001, 12'hF03} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hF05} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hF07} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hF08} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hF0C} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b001, 12'hF0F} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b001, 12'hF13} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hF14} : s_CHIP_26B_45133_reg = 8'h52;
         {3'b001, 12'hF18} : s_CHIP_26B_45133_reg = 8'hF2;
         {3'b001, 12'hF1B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hF1C} : s_CHIP_26B_45133_reg = 8'hF2;
         {3'b001, 12'hF1F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hF20} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b001, 12'hF23} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF24} : s_CHIP_26B_45133_reg = 8'h52;
         {3'b001, 12'hF27} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b001, 12'hF28} : s_CHIP_26B_45133_reg = 8'h52;
         {3'b001, 12'hF2B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b001, 12'hF2D} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b001, 12'hF2F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b001, 12'hF33} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hF34} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF37} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hF3B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hF3C} : s_CHIP_26B_45133_reg = 8'hF2;
         {3'b001, 12'hF3F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF40} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF42} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b001, 12'hF43} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF45} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hF47} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hF48} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF4A} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hF4B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF4C} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b001, 12'hF4F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b001, 12'hF51} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hF53} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hF54} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hF55} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hF57} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b001, 12'hF58} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF5B} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hF5C} : s_CHIP_26B_45133_reg = 8'hE1;
         {3'b001, 12'hF5F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF60} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hF61} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hF63} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hF64} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b001, 12'hF67} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'hF69} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b001, 12'hF6B} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b001, 12'hF6C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF6F} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b001, 12'hF70} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hF74} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hF78} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hF7C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hF80} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF82} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF83} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF84} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF86} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF87} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF88} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF8A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF8B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF8C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF8E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF8F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF90} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF92} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF93} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF94} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF96} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF97} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF98} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF9A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF9B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hF9C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hF9E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hF9F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hFA0} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hFA2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hFA3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hFA4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hFA6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hFA7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hFA8} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hFAA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hFAB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hFAC} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hFAE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hFAF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hFB0} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hFB2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hFB3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hFB4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hFB6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hFB7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hFB8} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hFBA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hFBB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hFBC} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b001, 12'hFBE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b001, 12'hFBF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b001, 12'hFC0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hFC3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'hFC4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hFC7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'hFC8} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hFCB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'hFCC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b001, 12'hFCF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'hFD0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hFD3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'hFD7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'hFD8} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b001, 12'hFDB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b001, 12'hFDC} : s_CHIP_26B_45133_reg = 8'hC4;
         {3'b001, 12'hFDF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b001, 12'hFE0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hFE4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hFE8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hFEC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hFF0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hFF4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hFF8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b001, 12'hFFC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b010, 12'h000} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h001} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h003} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b010, 12'h004} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h005} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h007} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h009} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h00A} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h00B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h00C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h00D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h00E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h00F} : s_CHIP_26B_45133_reg = 8'h42;
         {3'b010, 12'h011} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h012} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h013} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h015} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b010, 12'h017} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h018} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h019} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h01B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h01C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h01D} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b010, 12'h01F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h020} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h021} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h022} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h023} : s_CHIP_26B_45133_reg = 8'h42;
         {3'b010, 12'h025} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b010, 12'h026} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h027} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h028} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h029} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h02A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h02B} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b010, 12'h02C} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h02D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h02F} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h031} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h032} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h033} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h034} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h035} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h037} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h039} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h03A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h03B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h03D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h03F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b010, 12'h042} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h043} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h044} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h045} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h047} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b010, 12'h048} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h049} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h04B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h04D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h04F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h050} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b010, 12'h051} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h053} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h054} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h055} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h057} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h059} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h05A} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h05B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h05C} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b010, 12'h05D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h05F} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h061} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h062} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h063} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b010, 12'h065} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b010, 12'h067} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h068} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h069} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h06A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h06B} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b010, 12'h06C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h06D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h06F} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h071} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h073} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h075} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h077} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b010, 12'h079} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h07A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h07B} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h07D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h07E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h07F} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h081} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h082} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h083} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h085} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b010, 12'h086} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h087} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h089} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h08B} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b010, 12'h08C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h08D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h08E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h08F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h090} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h091} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h093} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h095} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h097} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b010, 12'h098} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b010, 12'h099} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h09B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h09C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b010, 12'h09D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h09E} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h09F} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b010, 12'h0A0} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h0A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h0A3} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h0A5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h0A6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h0A7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h0A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h0AB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b010, 12'h0AE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h0AF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h0B1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h0B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h0B4} : s_CHIP_26B_45133_reg = 8'h5B;
         {3'b010, 12'h0B5} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b010, 12'h0B6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h0B7} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b010, 12'h0B8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h0B9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h0BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h0BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h0BE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h0BF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h0C0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h0C1} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b010, 12'h0C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h0C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h0C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h0C6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h0C7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h0C9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h0CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h0CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h0CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h0CF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h0D0} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h0D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h0D3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h0D4} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b010, 12'h0D5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h0D6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h0D7} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b010, 12'h0D8} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h0D9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h0DA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h0DB} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b010, 12'h0DC} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h0DD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h0DE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h0DF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h0E1} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h0E3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b010, 12'h0E4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h0E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h0E7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h0E8} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h0E9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h0EB} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b010, 12'h0EC} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h0ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h0EF} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h0F0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h0F1} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b010, 12'h0F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h0F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h0F4} : s_CHIP_26B_45133_reg = 8'h58;
         {3'b010, 12'h0F5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h0F7} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h0F9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h0FA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h0FB} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h0FC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h0FD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h0FE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h0FF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h100} : s_CHIP_26B_45133_reg = 8'hC8;
         {3'b010, 12'h101} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h102} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h103} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h105} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h107} : s_CHIP_26B_45133_reg = 8'hB3;
         {3'b010, 12'h108} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h109} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h10B} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b010, 12'h10C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h10D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h10F} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h111} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h113} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h114} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h115} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h116} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h117} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b010, 12'h118} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h119} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h11B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h11D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h11E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h11F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h120} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h121} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h123} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h125} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h127} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h129} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h12B} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b010, 12'h12C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h12D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h12F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h131} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h132} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h133} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h134} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h135} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h137} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h138} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h139} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h13A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h13B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'h13D} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h13F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b010, 12'h140} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h141} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h143} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h144} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h145} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h147} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h148} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h149} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h14A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h14B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h14D} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b010, 12'h14F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h151} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h152} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h153} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h155} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h156} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h157} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h159} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h15B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h15C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h15D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h160} : s_CHIP_26B_45133_reg = 8'hFE;
         {3'b010, 12'h161} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h163} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b010, 12'h165} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b010, 12'h167} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h169} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h16A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h16B} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b010, 12'h16C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h16D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h16E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h16F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h171} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b010, 12'h173} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h175} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h177} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b010, 12'h178} : s_CHIP_26B_45133_reg = 8'hFE;
         {3'b010, 12'h179} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h17B} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b010, 12'h17C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h17D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h17F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h181} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h183} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b010, 12'h184} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h185} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b010, 12'h186} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h187} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h188} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h189} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b010, 12'h18A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h18B} : s_CHIP_26B_45133_reg = 8'h42;
         {3'b010, 12'h18C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h18D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h18E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h18F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h191} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h193} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h194} : s_CHIP_26B_45133_reg = 8'h98;
         {3'b010, 12'h195} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h196} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h197} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h199} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h19B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h19D} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b010, 12'h19E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h19F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h1A0} : s_CHIP_26B_45133_reg = 8'hC8;
         {3'b010, 12'h1A1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h1A3} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h1A5} : s_CHIP_26B_45133_reg = 8'h95;
         {3'b010, 12'h1A7} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b010, 12'h1A8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h1A9} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h1AA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h1AB} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b010, 12'h1AC} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h1AD} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b010, 12'h1AF} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h1B0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h1B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h1B2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h1B3} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b010, 12'h1B5} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b010, 12'h1B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h1B7} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'h1B8} : s_CHIP_26B_45133_reg = 8'h58;
         {3'b010, 12'h1BB} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b010, 12'h1BC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h1BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h1BF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h1C0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h1C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h1C3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h1C5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h1C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h1C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h1C9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h1CB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h1CC} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b010, 12'h1CD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h1CE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h1CF} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h1D0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h1D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h1D2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h1D3} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b010, 12'h1D5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h1D6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h1D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h1D8} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b010, 12'h1D9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h1DB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b010, 12'h1DC} : s_CHIP_26B_45133_reg = 8'h98;
         {3'b010, 12'h1DD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h1DF} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b010, 12'h1E1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h1E2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h1E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h1E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h1E7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h1E8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h1E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h1EB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h1EC} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b010, 12'h1ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h1EF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h1F0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h1F1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h1F2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h1F3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h1F4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h1F6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h1F7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h1F8} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h1F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h1FB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h1FC} : s_CHIP_26B_45133_reg = 8'h98;
         {3'b010, 12'h1FF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h202} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h203} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h204} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h205} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h207} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b010, 12'h209} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h20B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h20C} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h20D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h20F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h210} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'h211} : s_CHIP_26B_45133_reg = 8'h86;
         {3'b010, 12'h213} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h216} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h217} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h218} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h219} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h21B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h21C} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b010, 12'h21D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h21F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h220} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h221} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h223} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h224} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h227} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h228} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h229} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h22B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h22C} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b010, 12'h22D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h22F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h230} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h231} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h233} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h234} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h237} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h239} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h23B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h23C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h23D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h23F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h240} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h241} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h243} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h244} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h245} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h247} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h248} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h24B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h24C} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h24D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h24F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h250} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b010, 12'h251} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h253} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h254} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h255} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h257} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h258} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h25B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h25C} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h25D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h25F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h260} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b010, 12'h261} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h263} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h264} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h265} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h267} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h268} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h26B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h26D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h26F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h270} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h271} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h273} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h274} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h275} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h277} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h278} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h279} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h27B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h27C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h27F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h281} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h283} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h284} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h285} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h287} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h288} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b010, 12'h289} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h28B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h28C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h28D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h28F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h290} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h292} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h293} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h295} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h297} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h298} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h299} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h29B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h29C} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b010, 12'h29D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h29F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h2A0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2A1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h2A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2A4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2A6} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2A7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h2A9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h2AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h2AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2B0} : s_CHIP_26B_45133_reg = 8'h58;
         {3'b010, 12'h2B1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h2B3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h2B4} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b010, 12'h2B6} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2B7} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h2B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2BB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h2BC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2BD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h2BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2C3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h2C4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2C5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h2C6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h2C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2C8} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h2C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2CA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2CB} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'h2CC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h2CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2D1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h2D2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2D4} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h2D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2D7} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b010, 12'h2D8} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h2D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2DD} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h2DE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2E1} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h2E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2E7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h2E8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h2EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h2EF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h2F0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2F1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h2F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h2F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h2F4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2F5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h2F7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h2F8} : s_CHIP_26B_45133_reg = 8'h48;
         {3'b010, 12'h2F9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h2FA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h2FB} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'h2FC} : s_CHIP_26B_45133_reg = 8'h48;
         {3'b010, 12'h2FD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h2FF} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b010, 12'h301} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h303} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h304} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h305} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h309} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h30A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h30B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h30D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h30F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h311} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h313} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h314} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h315} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b010, 12'h316} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h317} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h318} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h319} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h31A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h31B} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h31C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h31D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h31F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h320} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h321} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h322} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h323} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h324} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h325} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h326} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h327} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h328} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h329} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h32A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h32B} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h32D} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h32E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h32F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h330} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h331} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h333} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h335} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h337} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b010, 12'h33B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b010, 12'h33C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h33D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h33F} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b010, 12'h340} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h341} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h342} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h343} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h346} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h347} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h348} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h349} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h34B} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b010, 12'h34C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h34D} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h34E} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b010, 12'h34F} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h352} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h353} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h354} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h355} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h357} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b010, 12'h358} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h359} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h35A} : s_CHIP_26B_45133_reg = 8'h4C;
         {3'b010, 12'h35B} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h35D} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h35E} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h35F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b010, 12'h362} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h363} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h364} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b010, 12'h365} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h366} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h367} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'h368} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h369} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b010, 12'h36B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h36E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h36F} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b010, 12'h371} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h372} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h373} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h374} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h375} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h377} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h378} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h379} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b010, 12'h37A} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b010, 12'h37B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b010, 12'h37D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h37F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h380} : s_CHIP_26B_45133_reg = 8'h58;
         {3'b010, 12'h381} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h383} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h384} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h385} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h387} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h388} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b010, 12'h389} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h38B} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b010, 12'h38C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h38D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h38F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h390} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h391} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h392} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h393} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b010, 12'h395} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h397} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b010, 12'h398} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h399} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h39B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h39C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h39E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h39F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h3A1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h3A3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h3A4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h3A5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h3A7} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b010, 12'h3A9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h3AA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h3AB} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b010, 12'h3AC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h3AD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h3AE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h3AF} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b010, 12'h3B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h3B2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h3B3} : s_CHIP_26B_45133_reg = 8'h29;
         {3'b010, 12'h3B5} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b010, 12'h3B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h3B8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h3B9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b010, 12'h3BA} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h3BB} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h3BD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h3BF} : s_CHIP_26B_45133_reg = 8'h38;
         {3'b010, 12'h3C0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h3C1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h3C3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b010, 12'h3C4} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h3C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h3C7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h3C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h3CA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h3CB} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b010, 12'h3CC} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h3CE} : s_CHIP_26B_45133_reg = 8'h8C;
         {3'b010, 12'h3CF} : s_CHIP_26B_45133_reg = 8'h6A;
         {3'b010, 12'h3D0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h3D1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h3D3} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b010, 12'h3D5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h3D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h3D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h3DB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h3DC} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h3DD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h3DE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h3DF} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b010, 12'h3E0} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b010, 12'h3E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h3E2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h3E3} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b010, 12'h3E4} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b010, 12'h3E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h3E6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h3E7} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b010, 12'h3E8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h3E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h3EA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h3EB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h3EC} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h3ED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h3EF} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h3F0} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h3F1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h3F3} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h3F4} : s_CHIP_26B_45133_reg = 8'hE8;
         {3'b010, 12'h3F5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h3F7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h3F8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h3FB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h3FC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h3FD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h3FF} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h401} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h403} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h404} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h405} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h406} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h407} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b010, 12'h409} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h40B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h40D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h40F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h410} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h413} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h414} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b010, 12'h415} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h417} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h419} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h41A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h41B} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h41C} : s_CHIP_26B_45133_reg = 8'hE9;
         {3'b010, 12'h41D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h41F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h420} : s_CHIP_26B_45133_reg = 8'h29;
         {3'b010, 12'h423} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h424} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h425} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h427} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h429} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h42B} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b010, 12'h42C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h42D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h42E} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b010, 12'h42F} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b010, 12'h430} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h431} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h433} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b010, 12'h434} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h435} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h437} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h438} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h439} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h43A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h43B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h43E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h43F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h441} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h443} : s_CHIP_26B_45133_reg = 8'h77;
         {3'b010, 12'h444} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h445} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h447} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b010, 12'h448} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h449} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h44B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h44D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h44E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h44F} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b010, 12'h450} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h451} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h452} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h453} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b010, 12'h454} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h455} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h456} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h457} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b010, 12'h459} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b010, 12'h45B} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b010, 12'h45C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h45D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b010, 12'h45E} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h45F} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h461} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h462} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h463} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h465} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h466} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h467} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b010, 12'h468} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h469} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h46B} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b010, 12'h46D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h46F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h470} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h471} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h473} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b010, 12'h474} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h475} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h477} : s_CHIP_26B_45133_reg = 8'h38;
         {3'b010, 12'h478} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h479} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h47B} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b010, 12'h47E} : s_CHIP_26B_45133_reg = 8'h4C;
         {3'b010, 12'h47F} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b010, 12'h482} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h483} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h484} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h485} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h487} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h488} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h489} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b010, 12'h48B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h48C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h48D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h48F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h490} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h491} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h493} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h494} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h495} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h497} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h498} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h499} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h49B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h49C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h49D} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h49F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h4A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4A3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b010, 12'h4A4} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h4A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4A7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h4A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4AB} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b010, 12'h4AC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h4AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4AF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h4B2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h4B3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b010, 12'h4B4} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h4B5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4B6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h4B7} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b010, 12'h4B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4BB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h4BD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h4BE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h4BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h4C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4C3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h4C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4C7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h4C8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h4C9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h4CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h4CB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h4CC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h4CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h4D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h4D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4D3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h4D4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h4D5} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h4D6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h4D7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h4D8} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'h4D9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h4DB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h4DC} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h4DD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4DE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h4DF} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b010, 12'h4E1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h4E2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h4E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h4E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4E7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h4E8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h4E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4EA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h4EB} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b010, 12'h4EC} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b010, 12'h4ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h4EE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h4EF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h4F0} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h4F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4F2} : s_CHIP_26B_45133_reg = 8'h48;
         {3'b010, 12'h4F3} : s_CHIP_26B_45133_reg = 8'hA8;
         {3'b010, 12'h4F4} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b010, 12'h4F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4F6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h4F7} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b010, 12'h4F8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h4F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h4FA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h4FB} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b010, 12'h4FD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h4FE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h4FF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h501} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h503} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h504} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h505} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h507} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h508} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h509} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h50A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h50B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h50C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h50D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h50F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h511} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h512} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h513} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h515} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h517} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h518} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h519} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h51A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h51B} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b010, 12'h51D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h51E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h51F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h521} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h523} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h524} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h525} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h526} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h527} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b010, 12'h528} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b010, 12'h529} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h52A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h52B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b010, 12'h52C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h52D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h52F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h530} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b010, 12'h531} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h532} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h533} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h534} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h535} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h538} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h539} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h53B} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b010, 12'h53C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h53D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h53F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h540} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b010, 12'h541} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h543} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b010, 12'h544} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h545} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h546} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h547} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h548} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'h549} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h54B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h54C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h54D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h54E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h54F} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b010, 12'h550} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h551} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h552} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h553} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h554} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h555} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h557} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h559} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h55A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h55B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'h55C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h55D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h55E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h55F} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b010, 12'h561} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h562} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h563} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'h564} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h565} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h567} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h568} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h569} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h56A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h56B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h56D} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b010, 12'h56F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h570} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b010, 12'h571} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h573} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b010, 12'h574} : s_CHIP_26B_45133_reg = 8'hF8;
         {3'b010, 12'h575} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h577} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b010, 12'h578} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h579} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h57B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'h57C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h57D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h57F} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b010, 12'h581} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h583} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b010, 12'h584} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h585} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b010, 12'h586} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h587} : s_CHIP_26B_45133_reg = 8'h42;
         {3'b010, 12'h588} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h589} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h58A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h58B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h58C} : s_CHIP_26B_45133_reg = 8'hFC;
         {3'b010, 12'h58D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h58F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h590} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h591} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b010, 12'h593} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h594} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h595} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b010, 12'h596} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h597} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h598} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h599} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h59A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h59B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h59C} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'h59D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h59F} : s_CHIP_26B_45133_reg = 8'hEE;
         {3'b010, 12'h5A0} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h5A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5A3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h5A5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h5A6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h5A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h5A9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h5AB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h5AC} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b010, 12'h5AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h5AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h5B0} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h5B1} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b010, 12'h5B2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h5B3} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b010, 12'h5B4} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h5B5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h5B7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h5B8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h5B9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h5BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h5BB} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'h5BC} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h5BF} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b010, 12'h5C0} : s_CHIP_26B_45133_reg = 8'h88;
         {3'b010, 12'h5C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5C3} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b010, 12'h5C4} : s_CHIP_26B_45133_reg = 8'hFC;
         {3'b010, 12'h5C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5C7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h5C8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h5C9} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b010, 12'h5CB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h5CC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h5CD} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b010, 12'h5CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h5D1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h5D2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h5D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h5D4} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b010, 12'h5D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5D7} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b010, 12'h5D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h5D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5DA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h5DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h5DD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h5DE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h5DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h5E0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h5E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5E2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h5E3} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'h5E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5E6} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h5E7} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h5E8} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h5E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5EB} : s_CHIP_26B_45133_reg = 8'hEE;
         {3'b010, 12'h5EC} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h5ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5EF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h5F0} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h5F1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h5F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h5F3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h5F4} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h5F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h5F6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b010, 12'h5F7} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b010, 12'h5F8} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h5F9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h5FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h5FB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h5FC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h5FD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h5FF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h601} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h602} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h603} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h605} : s_CHIP_26B_45133_reg = 8'h95;
         {3'b010, 12'h607} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h60B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b010, 12'h60C} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b010, 12'h60D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h60E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h60F} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'h610} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h611} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b010, 12'h613} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h615} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h617} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b010, 12'h61B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h61C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h61D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h61F} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h620} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h621} : s_CHIP_26B_45133_reg = 8'h55;
         {3'b010, 12'h622} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b010, 12'h623} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b010, 12'h625} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h627} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h628} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h629} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h62B} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h62C} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b010, 12'h62D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h62E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h62F} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'h630} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h631} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h633} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h634} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b010, 12'h635} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h637} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b010, 12'h638} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h639} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h63B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h63C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h63D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h63E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h63F} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b010, 12'h641} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h643} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b010, 12'h644} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b010, 12'h645} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h647} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h648} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h64A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h64B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h64C} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h64D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h64F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h650} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h651} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h652} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h653} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h654} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h655} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h657} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h659} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h65A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h65B} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b010, 12'h65E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h65F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h660} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h661} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h663} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h664} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h665} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h666} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b010, 12'h667} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h668} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h669} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h66B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h66D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h66E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h66F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h670} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h671} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h673} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h675} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h676} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h677} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h679} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h67B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h67C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h67D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h67E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h67F} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h680} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h681} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h683} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h684} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h685} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h686} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h687} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h688} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h689} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h68A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h68B} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h68C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h68D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h68F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h690} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h691} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h693} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h694} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h695} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h696} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h697} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h698} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h699} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h69A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h69B} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h69C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h69D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h69F} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h6A0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h6A1} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b010, 12'h6A2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h6A3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h6A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h6A6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h6A7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h6A8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h6A9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h6AA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h6AB} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h6AC} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h6AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h6AF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h6B0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h6B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h6B3} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h6B4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h6B5} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b010, 12'h6B6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h6B7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h6B9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h6BA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h6BB} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b010, 12'h6BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h6BE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h6BF} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h6C1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h6C2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h6C3} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b010, 12'h6C5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h6C7} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h6C8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h6C9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h6CB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h6CC} : s_CHIP_26B_45133_reg = 8'h29;
         {3'b010, 12'h6CF} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b010, 12'h6D0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h6D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h6D3} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b010, 12'h6D6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h6D7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h6D8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h6D9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h6DB} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h6DD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h6DF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h6E0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h6E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h6E3} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b010, 12'h6E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h6E7} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b010, 12'h6E8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b010, 12'h6E9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h6EB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h6EC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b010, 12'h6ED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h6EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h6F1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h6F2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h6F3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h6F4} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b010, 12'h6F5} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b010, 12'h6F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h6F8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h6F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h6FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h6FD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h6FE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h6FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h702} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h703} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h704} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h705} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h707} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h708} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h709} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h70A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h70B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h70C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h70D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h70F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h711} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h712} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h713} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h716} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h717} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h718} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b010, 12'h719} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h71B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h71D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h71E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h71F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'h720} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h721} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h723} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h724} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b010, 12'h725} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h727} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b010, 12'h729} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h72A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h72B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h72D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h72F} : s_CHIP_26B_45133_reg = 8'hB3;
         {3'b010, 12'h730} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h731} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h733} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h734} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b010, 12'h735} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h737} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b010, 12'h739} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h73A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h73B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h73D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h73F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h740} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b010, 12'h741} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h743} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h744} : s_CHIP_26B_45133_reg = 8'hC9;
         {3'b010, 12'h745} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h747} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b010, 12'h748} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b010, 12'h749} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h74B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h74D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h74E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h74F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h750} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h751} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h753} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h754} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h755} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h756} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h757} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h758} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h759} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h75B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h75D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h75E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h75F} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b010, 12'h762} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h763} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h764} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h765} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h767} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h768} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h769} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h76A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h76B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h76C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h76F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h771} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h772} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h773} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b010, 12'h775} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h776} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h777} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b010, 12'h779} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h77A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h77B} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b010, 12'h77D} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h77E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'h77F} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b010, 12'h780} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h781} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h783} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h784} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h785} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h787} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b010, 12'h788} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h789} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h78A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h78B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b010, 12'h78C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h78D} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b010, 12'h78F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'h790} : s_CHIP_26B_45133_reg = 8'hF8;
         {3'b010, 12'h791} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h793} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b010, 12'h794} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b010, 12'h795} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h797} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b010, 12'h798} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h799} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h79A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h79B} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h79D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h79F} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h7A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7A3} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h7A4} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b010, 12'h7A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7A7} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h7A8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b010, 12'h7A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7AB} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b010, 12'h7AC} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b010, 12'h7AD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h7AF} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b010, 12'h7B0} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b010, 12'h7B1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h7B2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h7B3} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b010, 12'h7B4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h7B5} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b010, 12'h7B7} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'h7B8} : s_CHIP_26B_45133_reg = 8'hFE;
         {3'b010, 12'h7B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7BB} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b010, 12'h7BC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h7BD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h7BF} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b010, 12'h7C0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h7C1} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b010, 12'h7C3} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'h7C4} : s_CHIP_26B_45133_reg = 8'hFE;
         {3'b010, 12'h7C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7C7} : s_CHIP_26B_45133_reg = 8'h8E;
         {3'b010, 12'h7C9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h7CB} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b010, 12'h7CC} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h7CD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h7CF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h7D0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h7D1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b010, 12'h7D2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h7D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h7D4} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h7D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7D7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h7D9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h7DA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h7DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h7DE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h7DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h7E0} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b010, 12'h7E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7E3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'h7E5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b010, 12'h7E6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h7E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h7E9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h7EB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'h7ED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b010, 12'h7EE} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b010, 12'h7EF} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b010, 12'h7F0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'h7F1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'h7F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h7F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7F6} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b010, 12'h7F7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'h7F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7FA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b010, 12'h7FB} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b010, 12'h7FC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b010, 12'h7FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h7FF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h801} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h802} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h803} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b010, 12'h804} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'h805} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b010, 12'h807} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h809} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h80A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h80B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h80D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b010, 12'h80F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h811} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'h812} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'h813} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'h814} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h818} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h81C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h820} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h824} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h828} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h82C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h830} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h834} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h838} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h83C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h840} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h844} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h848} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h84C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h850} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h854} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h858} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h85C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h860} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h864} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h868} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h86C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h870} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h874} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h878} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h87C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h880} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h884} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h888} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h88C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h890} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h894} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h898} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h89C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8A0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8A4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8A8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8AC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8B0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8B4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8B8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8BC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8C0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8C4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8C8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8CC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8D0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8D4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8D8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8DC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8E0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8E4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8E8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8EC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8F0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8F4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8F8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h8FC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h900} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h904} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h908} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h90C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h910} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h914} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h918} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h91C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h920} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h924} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h928} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h92C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h930} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h934} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h938} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h93C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h940} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h944} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h948} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h94C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h950} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h954} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h958} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h95C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h960} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h964} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h968} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h96C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h970} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h974} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h978} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h97C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h980} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h984} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h988} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h98C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h990} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h994} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h998} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h99C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9A0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9A4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9A8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9AC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9B0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9B4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9B8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9BC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9C0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9C4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9C8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9CC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9D0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9D4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9D8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9DC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9E0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9E4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9E8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9EC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9F0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9F4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9F8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'h9FC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA00} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA04} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA08} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA0C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA10} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA14} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA18} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA1C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA20} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA24} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA28} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA2C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA30} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA34} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA38} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA3C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA40} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA44} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA48} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA4C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA50} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA54} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA58} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA5C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA60} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA64} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA68} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA6C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA70} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA74} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA78} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA7C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA80} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA84} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA88} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA8C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA90} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA94} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA98} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hA9C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAA0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAA4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAA8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAAC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAB0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAB4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAB8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hABC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAC0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAC4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAC8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hACC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAD0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAD4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAD8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hADC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAE0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAE4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAE8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAEC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAF0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAF4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAF8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hAFC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB00} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB04} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB08} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB0C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB10} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB14} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB18} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB1C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB20} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB24} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB28} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB2C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB30} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB34} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB38} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB3C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB40} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB44} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB48} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB4C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB50} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB54} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB58} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB5C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB60} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB64} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB68} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB6C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB70} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB74} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB78} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB7C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB80} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB84} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB88} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB8C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB90} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB94} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB98} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hB9C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBA0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBA4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBA8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBAC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBB0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBB4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBB8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBBC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBC0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBC4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBC8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBCC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBD0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBD4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBD8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBDC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBE0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBE4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBE8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBEC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBF0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBF4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBF8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hBFC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b010, 12'hC00} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC04} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC08} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC0C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC10} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC14} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC18} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC1C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC20} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC24} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC28} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC2C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC30} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC34} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC38} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC3C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC40} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC44} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC48} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC4C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC50} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC54} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC58} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC5C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC60} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC64} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC68} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC6C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC70} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC74} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC78} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC7C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC80} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC84} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC88} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC8C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC90} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC94} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC98} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hC9C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCA0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCA4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCA8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCAC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCB0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCB4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCB8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCBC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCC0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCC4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCC8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCCC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCD0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCD4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCD8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCDC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCE0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCE4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCE8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCEC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCF0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCF4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCF8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hCFC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD00} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD04} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD08} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD0C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD10} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD14} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD18} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD1C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD20} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD24} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD28} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD2C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD30} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD34} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD38} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD3C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD40} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD44} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD48} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD4C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD50} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD54} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD58} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD5C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD60} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD64} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD68} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD6C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD70} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD74} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD78} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD7C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD80} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD84} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD88} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD8C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD90} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD94} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD98} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hD9C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDA0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDA4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDA8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDAC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDB0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDB4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDB8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDBC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDC0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDC4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDC8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDCC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDD0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDD4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDD8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDDC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDE0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDE4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDE8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDEC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDF0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDF4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDF8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hDFC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE00} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE04} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE08} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE0C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE10} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE14} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE18} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE1C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE20} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE24} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE28} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE2C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE30} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE34} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE38} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE3C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE40} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE44} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE48} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE4C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE50} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE54} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE58} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE5C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE60} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE64} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE68} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE6C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE70} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE74} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE78} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE7C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE80} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE84} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE88} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE8C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE90} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE94} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE98} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hE9C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hEA0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hEA4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hEA8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hEAC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hEB0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hEB4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hEB8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hEBC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b010, 12'hEC1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEC2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEC5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEC6} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEC9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hECA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hECD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hECE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hED1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hED2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hED5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hED6} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hED9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEDA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEDD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEDE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEE1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEE2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEE5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEE6} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEE9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEEA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEED} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEEE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEF1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEF2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEF5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEF6} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEF9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEFA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hEFD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hEFE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF00} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b010, 12'hF03} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b010, 12'hF04} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF07} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b010, 12'hF08} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF0C} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF0F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF10} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF13} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF14} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF17} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF18} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF1B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF1C} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF1F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF20} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b010, 12'hF22} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF23} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'hF24} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b010, 12'hF26} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF27} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'hF28} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b010, 12'hF2A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF2B} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'hF2C} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b010, 12'hF2E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF2F} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b010, 12'hF30} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b010, 12'hF33} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'hF34} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b010, 12'hF37} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'hF38} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b010, 12'hF3B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'hF3C} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b010, 12'hF3F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'hF40} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'hF41} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'hF42} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'hF43} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF44} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hF45} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'hF46} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'hF47} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'hF48} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF4B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF4C} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF4F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF50} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'hF51} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'hF52} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'hF53} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF54} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF57} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF59} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'hF5A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'hF5B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'hF5C} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF5F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF60} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'hF61} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'hF62} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'hF63} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF64} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b010, 12'hF65} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'hF66} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'hF67} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b010, 12'hF68} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF6B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF6C} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF6F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF70} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b010, 12'hF71} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'hF72} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'hF73} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF74} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF77} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF79} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b010, 12'hF7A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b010, 12'hF7B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b010, 12'hF7C} : s_CHIP_26B_45133_reg = 8'hA9;
         {3'b010, 12'hF7F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF80} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF83} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF84} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF87} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF88} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF8B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF8C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF8F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF90} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF93} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF94} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF97} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF98} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF9B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hF9C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hF9F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFA0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hFA3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFA7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFAB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFAF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFB3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFB7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFBB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFBF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFC0} : s_CHIP_26B_45133_reg = 8'hB8;
         {3'b010, 12'hFC3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'hFC4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hFC7} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b010, 12'hFC8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b010, 12'hFCB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFCC} : s_CHIP_26B_45133_reg = 8'hC8;
         {3'b010, 12'hFCF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'hFD0} : s_CHIP_26B_45133_reg = 8'hB8;
         {3'b010, 12'hFD3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b010, 12'hFD7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFDB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFDF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFE3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFE7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFEB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFEF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFF3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFF7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFFB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b010, 12'hFFF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h001} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h003} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h005} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h007} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h009} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h00B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h00D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h00F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h011} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h012} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h013} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h015} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h016} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h017} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h019} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h01A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h01B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h01D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h01E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h01F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h021} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h023} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h025} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h027} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h029} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h02B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h02D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h02F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h031} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h032} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h033} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h035} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h036} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h037} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h039} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h03A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h03B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h03D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h03E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h03F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h041} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h042} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h043} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h045} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h046} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h047} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h049} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h04A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h04B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h04D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h04E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h04F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h050} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h053} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h054} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h057} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h058} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h05B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h05C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h05F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h061} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h063} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h065} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h067} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h069} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h06B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h06D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h06F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h071} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h072} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h073} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h075} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h076} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h077} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h079} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h07A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h07B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h07D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h07E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h07F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h080} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h081} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h083} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h084} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h085} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h087} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h088} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h089} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h08B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h08C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h08D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h08F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h090} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h091} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h092} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h093} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h094} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h095} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h096} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h097} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h098} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h099} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h09A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h09B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h09C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h09D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h09E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h09F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h0A0} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0A3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0A4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0A7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0A8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0AB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0AC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0AF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0B0} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0B3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0B4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0B7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0B8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0BB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0BC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0BF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0C0} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0C3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h0C4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0C7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h0C8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0CB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h0CC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0CF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h0D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h0D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h0D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h0D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h0D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h0DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h0DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h0DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h0E0} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0E3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0E4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0E7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0E8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0EB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0EC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0EF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0F0} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0F3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0F4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0F7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0F8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0FB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h0FC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h0FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h0FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h0FF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h100} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h101} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h103} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h104} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h105} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h107} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h108} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h109} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h10B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h10C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h10D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h10F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h110} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h111} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h112} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h113} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h114} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h115} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h116} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h117} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h118} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h119} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h11A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h11B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h11C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h11D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h11E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h11F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h120} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h121} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h123} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h124} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h125} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h127} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h128} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h129} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h12B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h12C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h12D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h12F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h130} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h131} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h132} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h133} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h134} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h135} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h136} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h137} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h138} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h139} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h13A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h13B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h13C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h13D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h13E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h13F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h140} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h141} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h142} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h143} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h144} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h145} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h146} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h147} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h148} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h149} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h14A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h14B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h14C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h14D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h14E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h14F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h150} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h153} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h154} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h157} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h158} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h15B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h15C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h15F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h160} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h161} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h163} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h164} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h165} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h167} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h168} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h169} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h16B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h16C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h16D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h16F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h170} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h171} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h172} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h173} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h174} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h175} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h176} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h177} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h178} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h179} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h17A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h17B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h17C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h17D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h17E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h17F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h180} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h181} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h183} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h184} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h185} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h187} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h188} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h189} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h18B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h18C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h18D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h18F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h190} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h191} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h192} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h193} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h194} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h195} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h196} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h197} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h198} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h199} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h19A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h19B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h19C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h19D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h19E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h19F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h1A0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1A3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1A4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1A7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1A8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1AB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1AC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1AF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1B0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1B3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1B4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1B7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1B8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1BB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1BC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1BF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1C0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1C3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h1C4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1C7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h1C8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1CB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h1CC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1CF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h1D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h1D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h1D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h1DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h1E0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1E3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1E4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1E7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1E8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1EB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1EC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1EF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1F0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1F3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1F4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1F7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1F8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1FB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h1FC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h1FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h1FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h1FF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h200} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h201} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h203} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h204} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h205} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h207} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h208} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h209} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h20B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h20C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h20D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h20F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h210} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h211} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h212} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h213} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h214} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h215} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h216} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h217} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h218} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h219} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h21A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h21B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h21C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h21D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h21E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h21F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h220} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h221} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h223} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h224} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h225} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h227} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h228} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h229} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h22B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h22C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h22D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h22F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h230} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h231} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h232} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h233} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h234} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h235} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h236} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h237} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h238} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h239} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h23A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h23B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h23C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h23D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h23E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h23F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h240} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h241} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h242} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h243} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h244} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h245} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h246} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h247} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h248} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h249} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h24A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h24B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h24C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h24D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h24E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h24F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h250} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h253} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h254} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h257} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h258} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h25B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h25C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h25F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h260} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h261} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h263} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h264} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h265} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h267} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h268} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h269} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h26B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h26C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h26D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h26F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h270} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h271} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h272} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h273} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h274} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h275} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h276} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h277} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h278} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h279} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h27A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h27B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h27C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'h27D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h27E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h27F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h281} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h283} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h285} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h287} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h289} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h28B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h28D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h28F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h291} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h292} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h293} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h295} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h296} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h297} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h299} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h29A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h29B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h29D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h29E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h29F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h2D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h2D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h2DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h2DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h2FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h2FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h2FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h300} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h301} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h303} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h304} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h305} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h307} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h308} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h309} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h30B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h30C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h30D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h30F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h310} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h311} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h312} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h313} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h314} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h315} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h316} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h317} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h318} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h319} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h31A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h31B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h31C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h31D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h31E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h31F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h320} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h321} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h323} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h324} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h325} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h327} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h328} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h329} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h32B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h32C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h32D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h32F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h330} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h331} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h332} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h333} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h334} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h335} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h336} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h337} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h338} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h339} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h33A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h33B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h33C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h33D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h33E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h33F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h340} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h341} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h342} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h343} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h344} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h345} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h346} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h347} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h348} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h349} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h34A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h34B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h34C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h34D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h34E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h34F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'h350} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h353} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h354} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h357} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h358} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h35B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h35C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h35F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h360} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h361} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h363} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h364} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h365} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h367} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h368} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h369} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h36B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h36C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h36D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h36F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h370} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h371} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h372} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h373} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h374} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h375} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h376} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h377} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h378} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h379} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h37A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h37B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h37C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'h37D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h37E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h37F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'h381} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h383} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h385} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h387} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h389} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h38B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h38D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h38F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h391} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h392} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h393} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h395} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h396} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h397} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h399} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h39A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h39B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h39D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h39E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h39F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h3D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h3D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h3DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h3DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h3FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h3FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h3FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h401} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h403} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h405} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h407} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h409} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h40B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h40D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h40F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h411} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h412} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h413} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h415} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h416} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h417} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h419} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h41A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h41B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h41D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h41E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h41F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h421} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h423} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h425} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h427} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h429} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h42B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h42D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h42F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h431} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h432} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h433} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h435} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h436} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h437} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h439} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h43A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h43B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h43D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h43E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h43F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h441} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h442} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h443} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h445} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h446} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h447} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h449} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h44A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h44B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h44D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h44E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h44F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h450} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h453} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h454} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h457} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h458} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h45B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h45C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h45F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h461} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h463} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h465} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h467} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h469} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h46B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h46D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h46F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h471} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h472} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h473} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h475} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h476} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h477} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h479} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h47A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h47B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h47D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h47E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h47F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h481} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h483} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h485} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h487} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h489} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h48B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h48D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h48F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h491} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h492} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h493} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h495} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h496} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h497} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h499} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h49A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h49B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h49D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h49E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h49F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h4D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h4D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h4DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h4DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h4FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h4FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h4FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h501} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h503} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h505} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h507} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h509} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h50B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h50D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h50F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h511} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h512} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h513} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h515} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h516} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h517} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h519} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h51A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h51B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h51D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h51E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h51F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h521} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h523} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h525} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h527} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h529} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h52B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h52D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h52F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h531} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h532} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h533} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h535} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h536} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h537} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h539} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h53A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h53B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h53D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h53E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h53F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h541} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h542} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h543} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h545} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h546} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h547} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h549} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h54A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h54B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h54D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h54E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h54F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h550} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h553} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h554} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h557} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h558} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h55B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h55C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h55F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h561} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h563} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h565} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h567} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h569} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h56B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h56D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h56F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h571} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h572} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h573} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h575} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h576} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h577} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h579} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h57A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h57B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h57D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h57E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h57F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h581} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h583} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h585} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h587} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h589} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h58B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h58D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h58F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h591} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h592} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h593} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h595} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h596} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h597} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h599} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h59A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h59B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h59D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h59E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h59F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h5D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h5D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h5DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h5DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h5FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h5FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h5FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h601} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h603} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h605} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h607} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h609} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h60B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h60D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h60F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h611} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h612} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h613} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h615} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h616} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h617} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h619} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h61A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h61B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h61D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h61E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h61F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h621} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h623} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h625} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h627} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h629} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h62B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h62D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h62F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h631} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h632} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h633} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h635} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h636} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h637} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h639} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h63A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h63B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h63D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h63E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h63F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h641} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h642} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h643} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h645} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h646} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h647} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h649} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h64A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h64B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h64D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h64E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h64F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h650} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h653} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h654} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h657} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h658} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h65B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h65C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h65F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h661} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h663} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h665} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h667} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h669} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h66B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h66D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h66F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h671} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h672} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h673} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h675} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h676} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h677} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h679} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h67A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h67B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h67D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h67E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h67F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h681} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h683} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h685} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h687} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h689} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h68B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h68D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h68F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h691} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h692} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h693} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h695} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h696} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h697} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h699} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h69A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h69B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h69D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h69E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h69F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h6D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h6D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h6DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h6DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h6FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h6FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h6FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h701} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h703} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h705} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h707} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h709} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h70B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h70D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h70F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h711} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h712} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h713} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h715} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h716} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h717} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h719} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h71A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h71B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h71D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h71E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h71F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h721} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h723} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h725} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h727} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h729} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h72B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h72D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h72F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h731} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h732} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h733} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h735} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h736} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h737} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h739} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h73A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h73B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h73D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h73E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h73F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h741} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h742} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h743} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h745} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h746} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h747} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h749} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h74A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h74B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h74D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h74E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h74F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h750} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h753} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h754} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h757} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h758} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h75B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h75C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h75F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h761} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h763} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h765} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h767} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h769} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h76B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h76D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h76F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h771} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h772} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h773} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h775} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h776} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h777} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h779} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h77A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h77B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h77D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h77E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h77F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h781} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h783} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h785} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h787} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h789} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h78B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h78D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h78F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h791} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h792} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h793} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h795} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h796} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h797} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h799} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h79A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h79B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h79D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h79E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h79F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7A3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7AB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7C3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h7D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h7D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h7DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h7DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h7FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h7FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h7FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h800} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h801} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h803} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h804} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h805} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h807} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h808} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h809} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h80B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h80C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h80D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h80F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h810} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h811} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h812} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h813} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h814} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h815} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h816} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h817} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h818} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h819} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h81A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h81B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h81C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h81D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h81E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h81F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h821} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h823} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h825} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h827} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h829} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h82B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h82D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h82F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h831} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h832} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h833} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h835} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h836} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h837} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h839} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h83A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h83B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h83D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h83E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h83F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h840} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h841} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h842} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h843} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h844} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h845} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h846} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h847} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h848} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h849} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h84A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h84B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h84C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b011, 12'h84D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h84E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h84F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h850} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h853} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h854} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h857} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h858} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h85B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h85C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h85F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h861} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h863} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h865} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h867} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h869} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h86B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h86D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h86F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h871} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h872} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h873} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h875} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h876} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h877} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h879} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h87A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h87B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h87D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h87E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h87F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'h880} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h881} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h883} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h884} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h885} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h887} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h888} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h889} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h88B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h88C} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h88D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h88F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h890} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h891} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h892} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h893} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h894} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h895} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h896} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h897} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h898} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h899} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h89A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h89B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h89C} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h89D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h89E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h89F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8A0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8A3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8A4} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8A7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8A8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8AB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8AC} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8AF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8B0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8B3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8B4} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8B7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8B8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8BB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8BC} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8BF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8C0} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h8C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8C3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8C4} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h8C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8C7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8C8} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h8C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8CB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8CC} : s_CHIP_26B_45133_reg = 8'hF6;
         {3'b011, 12'h8CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8CF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h8D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h8D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h8D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h8D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h8DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h8DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h8DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h8E0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8E3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8E4} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8E7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8E8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8EB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8EC} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8EF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8F0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8F3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8F4} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8F7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8F8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8FB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h8FC} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b011, 12'h8FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h8FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h8FF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'h900} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h901} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h903} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h904} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h905} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h907} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h908} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h909} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h90B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h90C} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h90D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h90F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h910} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h911} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h912} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h913} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h914} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h915} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h916} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h917} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h918} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h919} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h91A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h91B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h91C} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h91D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h91E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h91F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h920} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h921} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h923} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h924} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h925} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h927} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h928} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h929} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h92B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h92C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h92D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h92F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h930} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h931} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h932} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h933} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h934} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h935} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h936} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h937} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h938} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h939} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h93A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h93B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h93C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h93D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h93E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h93F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h940} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h941} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h942} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h943} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h944} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h945} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h946} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h947} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h948} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h949} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h94A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h94B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h94C} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b011, 12'h94D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h94E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h94F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h950} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h953} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h954} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h957} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h958} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h95B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h95C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h95F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h960} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h961} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h963} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h964} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h965} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h967} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h968} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h969} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h96B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h96C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h96D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h96F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h970} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h971} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h972} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h973} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h974} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h975} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h976} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h977} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h978} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h979} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h97A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h97B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h97C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h97D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h97E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h97F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h980} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h981} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h983} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h984} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h985} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h987} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h988} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h989} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h98B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h98C} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h98D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h98F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h990} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h991} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h992} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h993} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h994} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h995} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h996} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h997} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h998} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h999} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h99A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h99B} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h99C} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h99D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h99E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h99F} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9A0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9A3} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9A4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9A7} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9A8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9A9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9AB} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9AC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9AF} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9B0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9B1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9B2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9B3} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9B4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9B5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9B7} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9B8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9B9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9BA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9BB} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9BC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9BD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9BE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9BF} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9C0} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h9C1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9C2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9C3} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9C4} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h9C5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9C6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9C7} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9C8} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h9C9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9CA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9CB} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9CC} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b011, 12'h9CD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9CE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9CF} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9D0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h9D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h9D4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h9D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h9D8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h9DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h9DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'h9DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'h9E0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9E1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9E3} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9E4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9E5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9E7} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9E8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9EB} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9EC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9EF} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9F0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9F1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9F2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9F3} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9F4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9F5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9F6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9F7} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9F8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9F9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9FB} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'h9FC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b011, 12'h9FD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'h9FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'h9FF} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b011, 12'hA00} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA01} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA03} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA04} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA05} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA07} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA08} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA09} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA0B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA0C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA0D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA0F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA10} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA11} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA12} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA13} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA14} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA15} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA16} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA17} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA18} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA19} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA1A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA1B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA1C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA1D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA1E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA1F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA21} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA23} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA25} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA27} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA29} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA2B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA2D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA2F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA31} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA32} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA33} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA35} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA36} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA37} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA39} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA3A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA3B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA3D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA3E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA3F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA40} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA41} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA42} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA43} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA44} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA45} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA46} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA47} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA48} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA49} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA4A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA4B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA4C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hA4D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA4E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA4F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA50} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hA53} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA54} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hA57} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA58} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hA5B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA5C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hA5F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA61} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA63} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA65} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA67} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA69} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA6B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA6D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA6F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA71} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA72} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA73} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA75} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA76} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA77} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA79} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA7A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA7B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA7D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA7E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA7F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hA81} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA82} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hA83} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA85} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA86} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hA87} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA89} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA8A} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hA8B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA8D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hA8E} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hA8F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA91} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA92} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hA93} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA95} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA96} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hA97} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA99} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA9A} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hA9B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hA9D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hA9E} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hA9F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAA1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAA3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAA5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAA7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAA9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAAB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAAD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAAF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAB1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hAB2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAB3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAB5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hAB6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAB7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAB9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hABA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hABB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hABD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hABE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hABF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAC1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hAC2} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hAC3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAC5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hAC6} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hAC7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAC9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hACA} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hACB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hACD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hACE} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hACF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAD0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hAD3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAD4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hAD7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAD8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hADB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hADC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hADF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAE1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAE3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAE5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAE7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAE9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAEB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAEF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAF1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hAF2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAF3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAF5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hAF6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAF7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAF9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hAFA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAFB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hAFD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hAFE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hAFF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hB00} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB01} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB02} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hB03} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB04} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB05} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB06} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hB07} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB08} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB09} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB0A} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hB0B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB0C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB0D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB0E} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hB0F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB10} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB11} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB12} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB13} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB14} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB15} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB16} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB17} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB18} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB19} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB1A} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB1B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB1C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB1D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB1E} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB1F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB20} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB21} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB22} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b011, 12'hB23} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB24} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB25} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB26} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b011, 12'hB27} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB28} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB29} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB2A} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b011, 12'hB2B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB2C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB2D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB2E} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b011, 12'hB2F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB30} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB31} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB32} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hB33} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB34} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB35} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB36} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hB37} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB38} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB39} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB3A} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hB3B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB3C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hB3D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB3E} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hB3F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB41} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB42} : s_CHIP_26B_45133_reg = 8'h47;
         {3'b011, 12'hB43} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b011, 12'hB45} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB46} : s_CHIP_26B_45133_reg = 8'h47;
         {3'b011, 12'hB47} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b011, 12'hB49} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB4A} : s_CHIP_26B_45133_reg = 8'h47;
         {3'b011, 12'hB4B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b011, 12'hB4D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB4E} : s_CHIP_26B_45133_reg = 8'h47;
         {3'b011, 12'hB4F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b011, 12'hB51} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB52} : s_CHIP_26B_45133_reg = 8'h43;
         {3'b011, 12'hB53} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b011, 12'hB55} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB56} : s_CHIP_26B_45133_reg = 8'h43;
         {3'b011, 12'hB57} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b011, 12'hB59} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB5A} : s_CHIP_26B_45133_reg = 8'h43;
         {3'b011, 12'hB5B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b011, 12'hB5D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB5E} : s_CHIP_26B_45133_reg = 8'h43;
         {3'b011, 12'hB5F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b011, 12'hB60} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hB61} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB62} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b011, 12'hB63} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB64} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hB65} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB66} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b011, 12'hB67} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB68} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hB69} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB6A} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b011, 12'hB6B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB6C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hB6D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB6E} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b011, 12'hB6F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB70} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hB71} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB72} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB73} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB74} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hB75} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB76} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB77} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB78} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hB79} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB7A} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB7B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB7C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hB7D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB7E} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB7F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hB80} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hB81} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB82} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB83} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hB84} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hB85} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB86} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB87} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hB88} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hB89} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB8A} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB8B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hB8C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hB8D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hB8E} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b011, 12'hB8F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hB90} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hB91} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hB92} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hB93} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hB94} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hB95} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hB96} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hB97} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hB98} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hB99} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hB9A} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hB9B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hB9C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hB9D} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hB9E} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hB9F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBA0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBA1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBA3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBA4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBA5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBA7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBA8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBA9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBAB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBAC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBAD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBAF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBB0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBB1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBB2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBB3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBB4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBB5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBB6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBB7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBB8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBB9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBBA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBBB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBBC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBBD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBBE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBBF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBC0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBC1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBC2} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hBC3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBC4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBC5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBC6} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hBC7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBC8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBC9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBCA} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hBCB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBCC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBCD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBCE} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b011, 12'hBCF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBD0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hBD3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBD4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hBD7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBD8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hBDB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBDC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hBDF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBE0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBE1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBE3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBE4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBE5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBE7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBE8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBE9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBEB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBEC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBEF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBF0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBF1} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBF2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBF3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBF4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBF5} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBF6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBF7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBF8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBF9} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBFA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBFB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hBFC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hBFD} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hBFE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b011, 12'hBFF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hC02} : s_CHIP_26B_45133_reg = 8'h4C;
         {3'b011, 12'hC03} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b011, 12'hC04} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'hC06} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hC07} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hC0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC0C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b011, 12'hC0F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC12} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b011, 12'hC13} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b011, 12'hC14} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hC17} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC18} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hC1B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC1C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b011, 12'hC1F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC22} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b011, 12'hC23} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b011, 12'hC27} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC28} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b011, 12'hC2B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC2F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC32} : s_CHIP_26B_45133_reg = 8'h4C;
         {3'b011, 12'hC33} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b011, 12'hC37} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC38} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hC3B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC3F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC42} : s_CHIP_26B_45133_reg = 8'h48;
         {3'b011, 12'hC43} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b011, 12'hC44} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b011, 12'hC47} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hC48} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b011, 12'hC4B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC4F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC52} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b011, 12'hC53} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b011, 12'hC57} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC58} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b011, 12'hC5A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b011, 12'hC5B} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b011, 12'hC5C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b011, 12'hC5F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hC62} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b011, 12'hC63} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b011, 12'hC64} : s_CHIP_26B_45133_reg = 8'hB8;
         {3'b011, 12'hC67} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b011, 12'hC68} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b011, 12'hC6B} : s_CHIP_26B_45133_reg = 8'hE6;
         {3'b011, 12'hC6C} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b011, 12'hC6F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b011, 12'hC72} : s_CHIP_26B_45133_reg = 8'h48;
         {3'b011, 12'hC73} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b011, 12'hC77} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC78} : s_CHIP_26B_45133_reg = 8'h68;
         {3'b011, 12'hC7B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b011, 12'hC7F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hC83} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b011, 12'hC87} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'hC8B} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b011, 12'hC8F} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b011, 12'hC92} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hC93} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hC96} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hC97} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b011, 12'hC9A} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hC9B} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b011, 12'hC9E} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hC9F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b011, 12'hCA2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCA3} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b011, 12'hCA6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCA7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hCAB} : s_CHIP_26B_45133_reg = 8'h7E;
         {3'b011, 12'hCAE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCAF} : s_CHIP_26B_45133_reg = 8'h7E;
         {3'b011, 12'hCB2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCB3} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b011, 12'hCB6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCB7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b011, 12'hCBB} : s_CHIP_26B_45133_reg = 8'h7E;
         {3'b011, 12'hCBE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCBF} : s_CHIP_26B_45133_reg = 8'h7E;
         {3'b011, 12'hCC2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCC3} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'hCC6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCC7} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hCCA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCCB} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b011, 12'hCCE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCCF} : s_CHIP_26B_45133_reg = 8'h6A;
         {3'b011, 12'hCD2} : s_CHIP_26B_45133_reg = 8'h4C;
         {3'b011, 12'hCD3} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'hCD6} : s_CHIP_26B_45133_reg = 8'h4C;
         {3'b011, 12'hCD7} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hCDA} : s_CHIP_26B_45133_reg = 8'h4C;
         {3'b011, 12'hCDB} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b011, 12'hCDE} : s_CHIP_26B_45133_reg = 8'h4C;
         {3'b011, 12'hCDF} : s_CHIP_26B_45133_reg = 8'h6A;
         {3'b011, 12'hCE2} : s_CHIP_26B_45133_reg = 8'h8C;
         {3'b011, 12'hCE3} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'hCE6} : s_CHIP_26B_45133_reg = 8'h8C;
         {3'b011, 12'hCE7} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hCEA} : s_CHIP_26B_45133_reg = 8'h8C;
         {3'b011, 12'hCEB} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b011, 12'hCEE} : s_CHIP_26B_45133_reg = 8'h8C;
         {3'b011, 12'hCEF} : s_CHIP_26B_45133_reg = 8'h6A;
         {3'b011, 12'hCF2} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCF3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hCF6} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCF7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hCFA} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCFB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hCFE} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b011, 12'hCFF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD00} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hD03} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD04} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b011, 12'hD07} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD08} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hD0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD0C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hD0F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD10} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hD13} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD17} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD1B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD1F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD20} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b011, 12'hD23} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD24} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b011, 12'hD27} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD28} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b011, 12'hD2B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD2C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b011, 12'hD2F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD30} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hD33} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD34} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hD37} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD38} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hD3B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD3C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b011, 12'hD3F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD40} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b011, 12'hD43} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hD44} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b011, 12'hD47} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hD48} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b011, 12'hD4B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hD4C} : s_CHIP_26B_45133_reg = 8'hE7;
         {3'b011, 12'hD4F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hD53} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD57} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD5B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD5F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD60} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b011, 12'hD63} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD64} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b011, 12'hD67} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD68} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b011, 12'hD6B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD6C} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b011, 12'hD6F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD70} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hD73} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD74} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hD77} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD7B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD7F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD83} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD87} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD8B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD8F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD93} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD97} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD9B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hD9F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDA3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDA7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDAB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDAF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDB3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDB7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDBB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDBF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDC3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDC7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDCB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDCF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDD3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDD7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDDB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDDF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDE3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDE7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDEB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDEF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDF3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDF7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDFB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hDFF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE00} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE03} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE04} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE07} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE08} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE0C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE0F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE10} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE13} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE14} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE17} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE18} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE1B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE1C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE1F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE20} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE23} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE24} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE27} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE28} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE2B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE2C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE2F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE30} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE33} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE34} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE37} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE38} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE3B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE3C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE3F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE40} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE43} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE44} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE47} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE48} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE4B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE4C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE4F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE50} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE53} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE54} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE57} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE58} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE5B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE5C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE5F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE60} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE63} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE64} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE67} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE68} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE6B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE6C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE6F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE70} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE73} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE74} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE77} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE78} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE7B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE7C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE7F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE80} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE83} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE84} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE87} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE88} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE8B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE8C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE8F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE90} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE93} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE94} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE97} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE98} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE9B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hE9C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hE9F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEA0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEA3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEA4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEA7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEA8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEAB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEAC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEAF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEB0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEB3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEB4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEB7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEB8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEBB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEBC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEBF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEC0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEC3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEC4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEC7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEC8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hECB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hECC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hECF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hED0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hED3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hED4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hED7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hED8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEDB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEDC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEDF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEE0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEE3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEE4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEE7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEE8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEEB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEEC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEEF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEF0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEF3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEF4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEF7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEF8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEFB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hEFC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b011, 12'hEFF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hF02} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF03} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF06} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF07} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF0A} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF0B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF0E} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF0F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF12} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF13} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF16} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF17} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF1A} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF1B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF1E} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF1F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF22} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF23} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF26} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF27} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF2A} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF2B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF2E} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF2F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF32} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF33} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF36} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF37} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF3A} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF3B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF3E} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF3F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b011, 12'hF40} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b011, 12'hF42} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF43} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF44} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b011, 12'hF46} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF47} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF48} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b011, 12'hF4A} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF4B} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF4C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b011, 12'hF4E} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF4F} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF50} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hF52} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF53} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF54} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hF56} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF57} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF58} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hF5A} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF5B} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF5C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b011, 12'hF5E} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF5F} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF60} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'hF62} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF63} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF64} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'hF66} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF67} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF68} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'hF6A} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF6B} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF6C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b011, 12'hF6E} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF6F} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF70} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hF72} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF73} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF74} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hF76} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF77} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF78} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hF7A} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF7B} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF7C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b011, 12'hF7E} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b011, 12'hF7F} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b011, 12'hF83} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hF87} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hF8B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hF8F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hF93} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hF97} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hF9B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hF9F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFA3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFA7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFAB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFAF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFB3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFB7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFBB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFBF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFC3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFC7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFCB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFCF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFD3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFD7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFDB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFDF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFE3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFE7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFEB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFEF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFF3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFF7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFFB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b011, 12'hFFF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1C0} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b100, 12'h1C3} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h1C4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h1C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1CA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h1CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1CC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b100, 12'h1CF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h1D0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'h1D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1D4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h1D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1D8} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h1DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1DC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b100, 12'h1DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1E0} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h1E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1E4} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'h1E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1E8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'h1EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1F0} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h1F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1F4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h1F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1F8} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h1FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h1FC} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h1FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h201} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h203} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h205} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h206} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h207} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b100, 12'h208} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h209} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h20B} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b100, 12'h20C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h20D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h20E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h20F} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b100, 12'h210} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h211} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h213} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h214} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h215} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h217} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b100, 12'h218} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h219} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h21B} : s_CHIP_26B_45133_reg = 8'hAC;
         {3'b100, 12'h21D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h21F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h220} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b100, 12'h221} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h223} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'h225} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h226} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h227} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'h228} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h229} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h22B} : s_CHIP_26B_45133_reg = 8'h7C;
         {3'b100, 12'h22C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h22D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h22E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h22F} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b100, 12'h230} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h231} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h233} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h234} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h235} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h237} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b100, 12'h238} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h239} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h23B} : s_CHIP_26B_45133_reg = 8'hAC;
         {3'b100, 12'h23D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h23F} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'h240} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h241} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h242} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h243} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'h244} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h245} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h247} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h248} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h249} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h24A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h24B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h24C} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h24D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h24F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h250} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h251} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h253} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h254} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h255} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h257} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h258} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h259} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h25B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h25C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h25D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h25F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h261} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h263} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h264} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h265} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h267} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h269} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h26B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h26D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h26F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h270} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h271} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h273} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h275} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h276} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h277} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h278} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h279} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h27A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h27B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h27C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h27D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h27E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'h27F} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b100, 12'h280} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'h281} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h285} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h287} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h288} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b100, 12'h289} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h28A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h28B} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h28C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'h28D} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h28F} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b100, 12'h290} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h291} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h292} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h293} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h294} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h295} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h297} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h299} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h29A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h29B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h29C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h29D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h29F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h2A1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h2A2} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'h2A3} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b100, 12'h2A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h2A6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h2A7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h2A8} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h2A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h2AA} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'h2AB} : s_CHIP_26B_45133_reg = 8'hFA;
         {3'b100, 12'h2AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h2AE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'h2AF} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b100, 12'h2B0} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h2B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h2B2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h2B3} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h2B4} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h2B5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h2B7} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h2B9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h2BA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h2BB} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h2BD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h2BF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h2C0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h2C1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h2C3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h2C5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h2C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h2C8} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h2C9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h2CA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h2CB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h2CC} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b100, 12'h2CD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h2CF} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h2D1} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h2D2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h2D3} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h2D4} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h2D5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h2D6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h2D7} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h2D8} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h2D9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h2DB} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h2DC} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h2DD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h2DF} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h2E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h2E2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h2E3} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b100, 12'h2E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h2E7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h2E8} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h2E9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h2EB} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h2EC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h2ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h2EF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h2F0} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h2F1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h2F3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h2F4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h2F5} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h2F6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h2F7} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b100, 12'h2F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h2FA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h2FB} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h2FD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h2FE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h2FF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h300} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h301} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h302} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h303} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h305} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h307} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h308} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h309} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h30B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h30C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h30D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h30F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h311} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h313} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h314} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h315} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h317} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h319} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h31B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h31D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h31F} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h321} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h323} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h325} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h327} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h328} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h329} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h32B} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h32C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h32D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h32F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h330} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h331} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h332} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h333} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h335} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h337} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h33A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h33B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h33C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h33D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h33F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h340} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h341} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h342} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h343} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b100, 12'h345} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h346} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h347} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h349} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h34A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h34B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h34C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h34D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h34E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h34F} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h350} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h351} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h353} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h355} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h357} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h358} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h359} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h35B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h35C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h35D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h35F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h361} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h363} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h364} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h365} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h367} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h368} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h369} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h36A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h36B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h36D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h36E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h36F} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b100, 12'h370} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h371} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h372} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h373} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h375} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h377} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h379} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h37B} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'h37F} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b100, 12'h381} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h382} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h383} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h384} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h385} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h387} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'h389} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h38B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h38C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h38D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h38E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h38F} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b100, 12'h391} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h392} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h393} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'h394} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h395} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h397} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b100, 12'h399} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h39B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h39C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h39D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h39E} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h39F} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'h3A0} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h3A1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h3A3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h3A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h3A7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h3A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h3AB} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b100, 12'h3AD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h3AF} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b100, 12'h3B0} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h3B1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h3B3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h3B4} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b100, 12'h3B5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h3B6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h3B7} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h3B8} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h3B9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h3BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h3BC} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b100, 12'h3BD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h3BE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h3BF} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h3C0} : s_CHIP_26B_45133_reg = 8'hD1;
         {3'b100, 12'h3C1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h3C2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h3C3} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b100, 12'h3C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h3C6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h3C7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h3C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h3CA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h3CB} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h3CC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h3CD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h3CF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h3D0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'h3D1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h3D2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h3D3} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'h3D4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h3D5} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b100, 12'h3D7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h3D9} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h3DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h3DD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h3DE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h3DF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h3E0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h3E1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h3E2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h3E3} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'h3E4} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h3E5} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b100, 12'h3E7} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h3E8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'h3E9} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h3EA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h3EB} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b100, 12'h3ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h3EE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h3EF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h3F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h3F2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h3F3} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h3F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h3F7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h3F8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h3F9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h3FA} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h3FB} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'h3FD} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b100, 12'h3FF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h401} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h403} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h405} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h406} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h407} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h408} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'h409} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h40A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h40B} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'h40D} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b100, 12'h40F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h410} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h411} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h413} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b100, 12'h414} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h415} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h417} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b100, 12'h418} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h419} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h41B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h41D} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h41E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h41F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h420} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h421} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h423} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h425} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h427} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h428} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h429} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h42B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h42C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h42D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h42E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h42F} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'h430} : s_CHIP_26B_45133_reg = 8'h91;
         {3'b100, 12'h431} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h432} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h433} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'h434} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h435} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h437} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'h438} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h439} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h43B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h43C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h43D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h43E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h43F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h440} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b100, 12'h441} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h443} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h445} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h447} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b100, 12'h449} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h44A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h44B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h44C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h44F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'h451} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h452} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h453} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'h454} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h455} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h457} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h458} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h45B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h45D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h45E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h45F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h461} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h462} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h463} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h465} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h467} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'h468} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h469} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h46B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h46D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h46F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h471} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h472} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h473} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h475} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h476} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h477} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h478} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h479} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h47B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'h47C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h47D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h47F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h480} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h481} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'h483} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'h485} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h487} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h488} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h489} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h48B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h48C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h48E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h48F} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h490} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h491} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h492} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h493} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h494} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h495} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h497} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'h499} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h49A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h49B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h49C} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h49D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h49F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h4A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4A3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h4A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4A6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h4A7} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h4A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4AB} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h4AC} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h4AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4AF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h4B1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h4B3} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b100, 12'h4B4} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h4B5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h4B6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h4B7} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'h4B8} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h4B9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h4BB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h4BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4BE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h4BF} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h4C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4C3} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h4C4} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h4C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4C7} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b100, 12'h4C8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h4C9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h4CB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h4CC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h4CD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h4CE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h4CF} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'h4D0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h4D1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h4D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h4D4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h4D5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h4D6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h4D7} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b100, 12'h4D8} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h4D9} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'h4DB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'h4DD} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h4DE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h4DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h4E0} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h4E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4E3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h4E4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h4E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4E7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h4E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4EA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h4EB} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h4ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4EF} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h4F0} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h4F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h4F3} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b100, 12'h4F4} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h4F5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h4F7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h4F8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h4F9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h4FA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h4FB} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'h4FC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h4FD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h4FF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h501} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h502} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h503} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h505} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h507} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h508} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h509} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h50B} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b100, 12'h50C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'h50D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h50F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h510} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h511} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h512} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h513} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'h514} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h515} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h517} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h518} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h519} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h51A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h51B} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b100, 12'h51C} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h51D} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'h51F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'h520} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h521} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h522} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h523} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h524} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h525} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h527} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h529} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h52B} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'h52D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h52F} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b100, 12'h530} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h531} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h533} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h535} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h536} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h537} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h538} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h539} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h53B} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'h53C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h53D} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h53F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h540} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h541} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h543} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h545} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h547} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h548} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h549} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h54B} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'h54C} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h54D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h54F} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h550} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b100, 12'h551} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h553} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h555} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h556} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h557} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h558} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h559} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h55B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h55C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h55D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h55F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h560} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h561} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h563} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h564} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h565} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h567} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h568} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h569} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h56B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h56C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h56D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h56F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h570} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b100, 12'h573} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h574} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h575} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h577} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h578} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h579} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h57B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h57C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h57D} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b100, 12'h57E} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b100, 12'h57F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h580} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h581} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h583} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h584} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'h585} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h587} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'h589} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h58B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h58D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h58E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h58F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h590} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h593} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b100, 12'h595} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h597} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'h599} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h59B} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b100, 12'h59C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h59D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h59F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h5A0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h5A1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h5A3} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h5A4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h5A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h5A8} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b100, 12'h5AA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5AB} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h5AC} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b100, 12'h5AD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h5AE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5AF} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h5B0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5B1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h5B2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5B3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h5B5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h5B6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h5B7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h5B8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h5B9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h5BA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5BB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h5BC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5BD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h5BF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h5C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h5C2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5C3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h5C4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h5C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h5C7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h5C8} : s_CHIP_26B_45133_reg = 8'hC1;
         {3'b100, 12'h5C9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h5CA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h5CB} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b100, 12'h5CC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h5CD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h5CF} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h5D0} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b100, 12'h5D1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h5D3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h5D4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h5D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h5D6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h5D8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5DB} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b100, 12'h5DC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h5DD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h5DF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h5E1} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h5E2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h5E3} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h5E7} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b100, 12'h5E9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h5EA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h5EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h5EC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h5ED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h5EE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h5EF} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'h5F0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h5F1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h5F3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h5F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h5F7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h5F8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h5F9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h5FA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h5FB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h5FC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h5FD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h5FF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h601} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h603} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b100, 12'h604} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h605} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h607} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h608} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h609} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h60B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h60D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h60F} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b100, 12'h611} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h613} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h614} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h615} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h617} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h618} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h619} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h61B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h61C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h61D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h61F} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b100, 12'h620} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h621} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h623} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b100, 12'h624} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h625} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h627} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h629} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h62A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h62B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h62D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h62F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h630} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h631} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b100, 12'h632} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h633} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'h635} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h637} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h639} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h63A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h63B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h63C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h63D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h63F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h641} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h643} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h645} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h647} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h648} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h649} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h64A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h64B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h64C} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h64D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h64F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h651} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h653} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'h655} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h657} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b100, 12'h658} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h659} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h65B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h65D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h65F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h661} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h663} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'h665} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h667} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b100, 12'h668} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h66B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h66C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h66D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h66E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h66F} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h671} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h673} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'h674} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h675} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h677} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'h678} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h679} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h67B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h67D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h67F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h680} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h681} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h682} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h683} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h684} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h685} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h687} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'h688} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h68B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h68C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h68D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h68E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h68F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h690} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b100, 12'h691} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h692} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h693} : s_CHIP_26B_45133_reg = 8'h7E;
         {3'b100, 12'h694} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'h695} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h697} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b100, 12'h699} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b100, 12'h69A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h69B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h69C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'h69D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h69E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h69F} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h6A0} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b100, 12'h6A1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h6A2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6A3} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h6A5} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h6A6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h6A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h6AB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h6AD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h6AE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h6AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h6B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h6B3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h6B4} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h6B5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h6B6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6B7} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h6B8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h6B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h6BB} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b100, 12'h6BC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h6BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h6BF} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h6C0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'h6C1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h6C2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h6C3} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h6C5} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h6C7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h6C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h6CA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h6CC} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h6CD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h6CF} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h6D0} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h6D1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h6D3} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h6D4} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h6D5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h6D6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6D7} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h6D8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6D9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h6DB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h6DC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'h6DD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h6DF} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'h6E0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6E3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h6E4} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h6E5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h6E6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6E7} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h6E8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h6EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h6EC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h6ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h6EF} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h6F0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6F3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h6F5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h6F7} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'h6F8} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h6FA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h6FB} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h6FC} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h6FD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h6FE} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h6FF} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'h700} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b100, 12'h701} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h703} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h705} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h707} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h709} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h70A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h70B} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'h70C} : s_CHIP_26B_45133_reg = 8'hA1;
         {3'b100, 12'h70D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h70F} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b100, 12'h711} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h713} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b100, 12'h714} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b100, 12'h715} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h716} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h717} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h718} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h719} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h71B} : s_CHIP_26B_45133_reg = 8'h18;
         {3'b100, 12'h71C} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h71F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h720} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b100, 12'h721} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h723} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h724} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h725} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h727} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h729} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h72B} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b100, 12'h72C} : s_CHIP_26B_45133_reg = 8'h52;
         {3'b100, 12'h72D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h72E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h72F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h730} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h731} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h733} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h734} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h735} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h737} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h738} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h739} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h73B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h73D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h73F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h741} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h743} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h744} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h745} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h746} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h747} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h748} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h749} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h74B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h74C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h74D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h74F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h750} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h751} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h752} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h753} : s_CHIP_26B_45133_reg = 8'h67;
         {3'b100, 12'h754} : s_CHIP_26B_45133_reg = 8'hC2;
         {3'b100, 12'h755} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h756} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h757} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'h758} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h759} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h75B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h75C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h75D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h75E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h75F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h761} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h763} : s_CHIP_26B_45133_reg = 8'h25;
         {3'b100, 12'h764} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h765} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h766} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h767} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h769} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h76B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'h76C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h76D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h76F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h770} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h771} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'h773} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h775} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h776} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h777} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b100, 12'h778} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b100, 12'h779} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h77B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h77C} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b100, 12'h77D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h77F} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h780} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h781} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h783} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b100, 12'h784} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h785} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h787} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h788} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b100, 12'h78A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h78B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h78D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h78E} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h78F} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'h790} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h791} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h793} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h794} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h795} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h797} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h799} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h79B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h79C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h79D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h79F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h7A0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'h7A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h7A3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'h7A4} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h7A5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h7A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h7A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h7AA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h7AB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h7AC} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'h7AF} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b100, 12'h7B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h7B3} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h7B4} : s_CHIP_26B_45133_reg = 8'hD1;
         {3'b100, 12'h7B5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h7B7} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h7B8} : s_CHIP_26B_45133_reg = 8'hF1;
         {3'b100, 12'h7B9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h7BB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h7BC} : s_CHIP_26B_45133_reg = 8'hC1;
         {3'b100, 12'h7BD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h7BF} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h7C0} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h7C1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h7C3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h7C4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h7C5} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'h7C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h7C8} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b100, 12'h7C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h7CB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h7CC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h7CF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h7D0} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b100, 12'h7D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h7D3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h7D4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h7D7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h7D8} : s_CHIP_26B_45133_reg = 8'h9A;
         {3'b100, 12'h7D9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h7DB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h7DC} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h7DF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h7E0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h7E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h7E3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h7E4} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h7E5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h7E6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h7E7} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h7E8} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b100, 12'h7E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h7EB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h7EC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h7ED} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h7EF} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h7F0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h7F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h7F2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h7F3} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h7F5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h7F7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h7F8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h7F9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h7FB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h7FC} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h7FF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h801} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h802} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h803} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'h804} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h805} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h806} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'h807} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b100, 12'h809} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h80B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h80C} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h80D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h80E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h80F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h811} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h813} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h814} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h815} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h817} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h818} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h819} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h81A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h81B} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h81D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h81E} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h81F} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'h820} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'h821} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h823} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h825} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h827} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h828} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h829} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'h82A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h82B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h82D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h82E} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h82F} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'h830} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b100, 12'h831} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h833} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h834} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h835} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h837} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'h838} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b100, 12'h839} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h83B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h83C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h83D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h83F} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'h840} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'h841} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h843} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h844} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h845} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h847} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h848} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h84B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h84C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h84D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h84F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h850} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h851} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h852} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h853} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h854} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'h856} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h857} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h859} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h85A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h85B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h85C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h85D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h85F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'h861} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h862} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h863} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h864} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h865} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h866} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h867} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h868} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'h869} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h86B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h86C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h86F} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b100, 12'h871} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h873} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h875} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h876} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h877} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'h879} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h87B} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b100, 12'h87C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h87D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h87F} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b100, 12'h880} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h881} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h883} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h884} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h885} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h887} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h888} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h889} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h88A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h88B} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h88C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h88D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h88E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h88F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h890} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h891} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h893} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h894} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h895} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h896} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h897} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h898} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h899} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h89B} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'h89D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h89F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h8A0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h8A1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h8A3} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'h8A4} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'h8A5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h8A7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h8A8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h8A9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h8AB} : s_CHIP_26B_45133_reg = 8'h37;
         {3'b100, 12'h8AC} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'h8AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h8AF} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'h8B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h8B3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h8B4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h8B5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h8B7} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'h8B8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h8B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h8BB} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'h8BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h8BF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h8C1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h8C2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h8C3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h8C5} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h8C7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h8C8} : s_CHIP_26B_45133_reg = 8'h21;
         {3'b100, 12'h8CB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h8CC} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h8CD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h8CE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h8CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h8D0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h8D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h8D3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h8D4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h8D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h8D7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h8D9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h8DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h8DD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h8DF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h8E0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h8E1} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h8E2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h8E3} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h8E4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h8E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h8E7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h8E8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h8E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h8EB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h8EC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h8ED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h8EE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h8EF} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h8F0} : s_CHIP_26B_45133_reg = 8'hC2;
         {3'b100, 12'h8F1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h8F2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h8F3} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'h8F5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h8F6} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h8F7} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'h8F8} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h8F9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h8FA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h8FB} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h8FD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h8FF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h900} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h901} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h903} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h905} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h907} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'h908} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h909} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h90B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h90C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h90D} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'h90F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h910} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h911} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h913} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h914} : s_CHIP_26B_45133_reg = 8'h82;
         {3'b100, 12'h915} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h916} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h917} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'h919} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h91A} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h91B} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'h91C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h91D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h91F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'h920} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h921} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h922} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h923} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h925} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h927} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h928} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h929} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h92B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h92C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h92D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h92E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h92F} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h931} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h932} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h933} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'h934} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'h935} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'h937} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h939} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h93B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'h93C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h93D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h93F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h940} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'h943} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'h945} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h947} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h948} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h949} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h94B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h94C} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'h94D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h94F} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'h950} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h951} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h953} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h955} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h956} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h957} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'h958} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h959} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h95B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h95C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h95D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h95F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h960} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h961} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h963} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b100, 12'h964} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h965} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b100, 12'h966} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b100, 12'h967} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h969} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h96B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h96C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h96D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h96F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h970} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h971} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h972} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h973} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h975} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h977} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'h978} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h979} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h97B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h97C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h97D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h97F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h980} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'h981} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h983} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h984} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h985} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h987} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h988} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h989} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h98B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h98C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h98D} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b100, 12'h98E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h98F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h991} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h993} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b100, 12'h994} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h995} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h997} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h999} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h99B} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b100, 12'h99D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h99F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'h9A0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'h9A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h9A3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'h9A5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h9A6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h9A7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h9A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h9AB} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h9AC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h9AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h9AF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'h9B0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h9B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h9B3} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h9B4} : s_CHIP_26B_45133_reg = 8'h52;
         {3'b100, 12'h9B5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h9B7} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b100, 12'h9B8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h9B9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'h9BB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'h9BC} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h9BD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h9BE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h9BF} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b100, 12'h9C0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'h9C1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h9C3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'h9C4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'h9C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h9C7} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'h9C8} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h9C9} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h9CB} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h9CD} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'h9CE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'h9CF} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b100, 12'h9D0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'h9D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h9D2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h9D3} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'h9D4} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h9D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h9D7} : s_CHIP_26B_45133_reg = 8'h78;
         {3'b100, 12'h9D8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'h9D9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h9DA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h9DB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'h9DC} : s_CHIP_26B_45133_reg = 8'hB2;
         {3'b100, 12'h9DD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h9DF} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'h9E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h9E2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'h9E3} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b100, 12'h9E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'h9E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h9E8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h9E9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h9EB} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'h9EC} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'h9ED} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'h9EE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h9EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'h9F0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'h9F1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'h9F2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h9F3} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b100, 12'h9F4} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'h9F5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'h9F6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h9F7} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h9F8} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'h9FA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'h9FB} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'h9FC} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'h9FD} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'h9FF} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b100, 12'hA01} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA02} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hA03} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hA05} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hA06} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hA07} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hA08} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hA09} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hA0A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hA0B} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hA0D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hA0F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hA11} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA13} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hA14} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hA15} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hA17} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hA19} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA1B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hA1D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA1F} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hA21} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hA23} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hA24} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'hA25} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hA26} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hA27} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hA28} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hA29} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA2B} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hA2C} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hA2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA2F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hA30} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b100, 12'hA31} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hA33} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b100, 12'hA34} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hA36} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hA37} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hA39} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA3B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hA3C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hA3D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hA3F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hA41} : s_CHIP_26B_45133_reg = 8'hB4;
         {3'b100, 12'hA43} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hA45} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hA47} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'hA48} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hA49} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hA4A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hA4B} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b100, 12'hA4D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hA4F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hA50} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hA52} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hA53} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'hA54} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hA55} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hA56} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hA57} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hA58} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hA59} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hA5B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hA5D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA5F} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'hA60} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hA62} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hA63} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b100, 12'hA65} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA66} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hA67} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'hA68} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'hA69} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA6B} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hA6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA6F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hA70} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hA71} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'hA73} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hA74} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hA75} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hA76} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hA77} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hA78} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'hA79} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hA7A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hA7B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hA7C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hA7D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA7E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'hA7F} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b100, 12'hA81} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hA82} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'hA83} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b100, 12'hA85} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hA87} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hA89} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA8B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hA8D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hA8F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'hA90} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hA91} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hA93} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'hA94} : s_CHIP_26B_45133_reg = 8'hC2;
         {3'b100, 12'hA95} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hA97} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hA99} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA9B} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hA9D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hA9E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'hA9F} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b100, 12'hAA1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hAA3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hAA5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hAA6} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'hAA7} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b100, 12'hAA8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hAA9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hAAA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hAAB} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b100, 12'hAAC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hAAD} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hAAE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hAAF} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hAB1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hAB3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hAB5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hAB7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hAB9} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hABB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hABD} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hABE} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'hABF} : s_CHIP_26B_45133_reg = 8'hD9;
         {3'b100, 12'hAC0} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hAC1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hAC3} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b100, 12'hAC4} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'hAC5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hAC7} : s_CHIP_26B_45133_reg = 8'h2C;
         {3'b100, 12'hAC9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hACB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hACD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hACF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hAD0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hAD1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hAD2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hAD3} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b100, 12'hAD5} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hAD7} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'hAD9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hADB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hADC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hADD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hADF} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hAE0} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hAE1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hAE2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hAE3} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hAE4} : s_CHIP_26B_45133_reg = 8'hA3;
         {3'b100, 12'hAE5} : s_CHIP_26B_45133_reg = 8'hB4;
         {3'b100, 12'hAE7} : s_CHIP_26B_45133_reg = 8'h7D;
         {3'b100, 12'hAE9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hAEB} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'hAEC} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hAED} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hAEE} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hAEF} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'hAF0} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hAF1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hAF2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hAF3} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b100, 12'hAF4} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hAF5} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'hAF7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hAF9} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hAFA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hAFB} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'hAFC} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hAFD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hAFE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hAFF} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hB00} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hB01} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hB03} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hB05} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB06} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hB07} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'hB09} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hB0B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hB0C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hB0D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB0E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hB0F} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hB10} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hB11} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB13} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b100, 12'hB15} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hB17} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hB19} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB1A} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB1B} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'hB1C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hB1D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hB1F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hB20} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hB21} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB23} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hB24} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hB25} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB27} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'hB28} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hB29} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB2B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hB2C} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b100, 12'hB2D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hB2E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hB2F} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hB30} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'hB32} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hB33} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hB35} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB36} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hB37} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hB38} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hB39} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hB3A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hB3B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hB3C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hB3D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hB3E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hB3F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hB40} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hB43} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'hB45} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB47} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hB48} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'hB49} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB4A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hB4B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hB4C} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hB4D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hB4F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hB51} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB52} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hB53} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b100, 12'hB54} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hB57} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b100, 12'hB58} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'hB59} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB5B} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hB5D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB5F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hB61} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB62} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hB63} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'hB64} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hB65} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB67} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'hB69} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB6B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hB6C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hB6D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hB6F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hB70} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'hB71} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB72} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hB73} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'hB74} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b100, 12'hB75} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hB76} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hB77} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hB79} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hB7B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hB7D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hB7E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hB7F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hB80} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hB81} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB82} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hB83} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b100, 12'hB84} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hB85} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b100, 12'hB87} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hB88} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'hB89} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB8B} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hB8D} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hB8E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hB8F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'hB90} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hB93} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hB95} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'hB96} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB97} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hB98} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hB99} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hB9B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'hB9C} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'hB9D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hB9F} : s_CHIP_26B_45133_reg = 8'h37;
         {3'b100, 12'hBA0} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'hBA1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hBA3} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hBA5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBA7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hBA8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hBA9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBAB} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hBAC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hBAD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBAF} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'hBB0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'hBB1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBB2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hBB3} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hBB5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hBB6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hBB7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hBB9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hBBB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hBBC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hBBD} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hBBF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hBC0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hBC1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hBC3} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b100, 12'hBC4} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'hBC5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hBC6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hBC7} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hBC9} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hBCA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hBCB} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hBCD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBCF} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b100, 12'hBD1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hBD2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hBD3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hBD4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'hBD5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hBD6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hBD7} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'hBD9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hBDB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hBDC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hBDD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hBDF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hBE1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hBE3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hBE4} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hBE5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBE7} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'hBE9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBEA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hBEB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hBED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBEE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hBEF} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hBF1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBF3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hBF5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hBF7} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hBF8} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'hBF9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hBFA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hBFB} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hBFC} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hBFD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hBFE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hBFF} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b100, 12'hC01} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC02} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hC03} : s_CHIP_26B_45133_reg = 8'h69;
         {3'b100, 12'hC04} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hC05} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC07} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'hC08} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hC09} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC0A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hC0B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hC0C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hC0D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hC0E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hC0F} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hC10} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hC11} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hC12} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hC13} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hC14} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hC15} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC16} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'hC17} : s_CHIP_26B_45133_reg = 8'hBA;
         {3'b100, 12'hC19} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC1A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'hC1B} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b100, 12'hC1C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'hC1D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC1E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hC1F} : s_CHIP_26B_45133_reg = 8'h64;
         {3'b100, 12'hC21} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b100, 12'hC23} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hC25} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC27} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hC29} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hC2B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'hC2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC2E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hC2F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hC31} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC33} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'hC34} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hC35} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hC37} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'hC38} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hC39} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hC3B} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hC3D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC3E} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'hC3F} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b100, 12'hC40} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hC41} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC43} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hC45} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC47} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hC49} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hC4B} : s_CHIP_26B_45133_reg = 8'hE5;
         {3'b100, 12'hC4D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC4F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hC50} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hC51} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC53} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b100, 12'hC55} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b100, 12'hC57} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'hC59} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hC5A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b100, 12'hC5B} : s_CHIP_26B_45133_reg = 8'h99;
         {3'b100, 12'hC5D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC5F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hC60} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'hC61} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC63} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b100, 12'hC65} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC67} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hC69} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hC6B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hC6C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hC6D} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'hC6F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hC70} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hC71} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hC72} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hC73} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b100, 12'hC74} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hC75} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hC77} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hC78} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'hC79} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hC7B} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b100, 12'hC7D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC7F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hC81} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC83} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hC85} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hC87} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hC88} : s_CHIP_26B_45133_reg = 8'hA3;
         {3'b100, 12'hC89} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'hC8B} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'hC8C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC8D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hC8E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hC8F} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hC90} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hC91} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hC93} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hC94} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hC95} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC96} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hC97} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hC99} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hC9B} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hC9C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hC9D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hC9F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hCA0} : s_CHIP_26B_45133_reg = 8'hA3;
         {3'b100, 12'hCA1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hCA3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hCA4} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hCA5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hCA6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hCA7} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b100, 12'hCA8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hCA9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hCAB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hCAD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hCAF} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'hCB0} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b100, 12'hCB1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hCB2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hCB3} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hCB4} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hCB5} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'hCB7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hCB8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hCB9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hCBB} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'hCBC} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hCBD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hCBF} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hCC0} : s_CHIP_26B_45133_reg = 8'hB2;
         {3'b100, 12'hCC1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hCC3} : s_CHIP_26B_45133_reg = 8'h7E;
         {3'b100, 12'hCC4} : s_CHIP_26B_45133_reg = 8'hD3;
         {3'b100, 12'hCC7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hCC8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'hCC9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hCCA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hCCB} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hCCC} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b100, 12'hCCD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hCCF} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hCD1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hCD3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hCD5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hCD6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hCD7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hCD8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'hCD9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hCDB} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hCDD} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hCDF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hCE1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hCE3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hCE4} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hCE7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hCE8} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'hCE9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hCEA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hCEB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hCEC} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hCED} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hCEF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hCF1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hCF3} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'hCF5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hCF7} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b100, 12'hCF8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hCF9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hCFA} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hCFB} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hCFC} : s_CHIP_26B_45133_reg = 8'h42;
         {3'b100, 12'hCFD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hCFF} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'hD00} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'hD01} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD03} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hD04} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hD05} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hD07} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hD08} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hD09} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD0A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hD0B} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hD0D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD0F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hD11} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hD12} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hD13} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'hD14} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b100, 12'hD15} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hD17} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hD18} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hD19} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hD1B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hD1C} : s_CHIP_26B_45133_reg = 8'hD3;
         {3'b100, 12'hD1D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hD1F} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hD21} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hD23} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hD24} : s_CHIP_26B_45133_reg = 8'hD2;
         {3'b100, 12'hD25} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hD27} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hD28} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hD29} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hD2B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hD2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD2F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hD31} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hD33} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hD35} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hD37} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hD38} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hD39} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hD3A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hD3B} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hD3D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD3F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hD41} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hD42} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hD43} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'hD44} : s_CHIP_26B_45133_reg = 8'h92;
         {3'b100, 12'hD45} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hD47} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hD48} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b100, 12'hD4B} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'hD4C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'hD4D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD4F} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'hD50} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'hD51} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD53} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hD54} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b100, 12'hD55} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD57} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hD58} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hD59} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hD5A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hD5B} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hD5C} : s_CHIP_26B_45133_reg = 8'hC2;
         {3'b100, 12'hD5D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hD5F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b100, 12'hD60} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'hD61} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD63} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hD64} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hD65} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hD67} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hD68} : s_CHIP_26B_45133_reg = 8'hD3;
         {3'b100, 12'hD6A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hD6B} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hD6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD6F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hD70} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hD71} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hD73} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b100, 12'hD74} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hD75} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hD77} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b100, 12'hD78} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hD79} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hD7B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hD7D} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hD7E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hD7F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'hD80} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hD81} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD83} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hD84} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b100, 12'hD87} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hD88} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hD89} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD8B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hD8C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hD8D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD8F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hD90} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'hD91} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD93} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hD94} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hD95} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hD97} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hD98} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hD99} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hD9B} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b100, 12'hD9C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hD9D} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b100, 12'hD9E} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b100, 12'hD9F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hDA1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hDA3} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hDA4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b100, 12'hDA5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDA7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hDA8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hDA9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hDAA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hDAB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hDAD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDAF} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'hDB0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hDB1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDB2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hDB3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hDB4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hDB5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDB7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hDB8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'hDB9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDBB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hDBC} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hDBD} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b100, 12'hDBE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hDBF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hDC1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDC3} : s_CHIP_26B_45133_reg = 8'h5E;
         {3'b100, 12'hDC5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDC7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hDC8} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b100, 12'hDC9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDCB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hDCD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hDCE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hDCF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hDD1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDD3} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hDD4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hDD5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDD7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hDD8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hDD9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDDB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hDDD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDDF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hDE0} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hDE1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hDE3} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b100, 12'hDE4} : s_CHIP_26B_45133_reg = 8'h53;
         {3'b100, 12'hDE5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hDE7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hDE8} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hDE9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDEB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hDED} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hDEF} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hDF1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDF3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hDF4} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'hDF5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hDF7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hDF8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hDFB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hDFC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hDFD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hDFF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hE00} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b100, 12'hE01} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hE02} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hE03} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b100, 12'hE05} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE07} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b100, 12'hE09} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hE0A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hE0B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hE0C} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'hE0D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hE0E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hE0F} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b100, 12'hE11} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hE13} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hE15} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE17} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hE18} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hE19} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hE1B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hE1C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hE1D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hE1F} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hE21} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE23} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hE24} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hE25} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE27} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'hE29} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hE2B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hE2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE2F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hE30} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b100, 12'hE31} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hE32} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hE33} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hE34} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hE35} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hE37} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hE39} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE3A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hE3B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hE3C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hE3D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE3E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hE3F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hE41} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE43} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hE44} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b100, 12'hE45} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE47} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hE49} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE4B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hE4C} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hE4D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hE4F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hE50} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hE51} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE53} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hE54} : s_CHIP_26B_45133_reg = 8'hC3;
         {3'b100, 12'hE55} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hE57} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hE58} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hE59} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hE5B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hE5C} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hE5D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hE5E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hE5F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hE60} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hE61} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hE63} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hE64} : s_CHIP_26B_45133_reg = 8'h93;
         {3'b100, 12'hE65} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hE67} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hE69} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE6A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hE6B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'hE6D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hE6E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hE6F} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b100, 12'hE70} : s_CHIP_26B_45133_reg = 8'h93;
         {3'b100, 12'hE71} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hE72} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hE73} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b100, 12'hE75} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE76} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hE77} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b100, 12'hE78} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hE79} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hE7A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hE7B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'hE7D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE7F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hE81} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hE82} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hE83} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b100, 12'hE84} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hE85} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hE86} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hE87} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hE89} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE8A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hE8B} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b100, 12'hE8C} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hE8D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hE8E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hE8F} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b100, 12'hE90} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hE92} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hE93} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b100, 12'hE95} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE96} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hE97} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b100, 12'hE98} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hE9B} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b100, 12'hE9C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hE9D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hE9E} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hE9F} : s_CHIP_26B_45133_reg = 8'h2B;
         {3'b100, 12'hEA0} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'hEA1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hEA2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hEA3} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b100, 12'hEA4} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hEA5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hEA6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hEA7} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b100, 12'hEA8} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b100, 12'hEA9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hEAA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hEAB} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hEAC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hEAD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hEAF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hEB1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hEB3} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hEB4} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hEB7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hEB8} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b100, 12'hEB9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hEBB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hEBC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hEBD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hEBF} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hEC0} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'hEC1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hEC2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hEC3} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b100, 12'hEC4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hEC5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hEC7} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hEC8} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hEC9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hECB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hECD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hECE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hECF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hED1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hED3} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'hED5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hED7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hED9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hEDB} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hEDC} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hEDF} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'hEE0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hEE1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hEE3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'hEE4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hEE5} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hEE6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hEE7} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b100, 12'hEE9} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b100, 12'hEEB} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b100, 12'hEEC} : s_CHIP_26B_45133_reg = 8'hF3;
         {3'b100, 12'hEEF} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b100, 12'hEF1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hEF3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hEF4} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'hEF6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hEF7} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b100, 12'hEF8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hEF9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hEFB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hEFC} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hEFD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hEFF} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hF00} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b100, 12'hF02} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF03} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hF05} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF06} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF07} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hF09} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF0B} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hF0C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hF0D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF0F} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b100, 12'hF11} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF13} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hF15} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF17} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b100, 12'hF18} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b100, 12'hF19} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hF1B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b100, 12'hF1C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hF1D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hF1F} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hF21} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF23} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hF25} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF27} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hF28} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hF29} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hF2A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hF2B} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b100, 12'hF2D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF2E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hF2F} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b100, 12'hF30} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hF31} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hF32} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF33} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hF35} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF36} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hF37} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b100, 12'hF38} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hF39} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hF3A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hF3B} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b100, 12'hF3C} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hF3D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hF3E} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hF3F} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b100, 12'hF40} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hF41} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hF43} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hF44} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hF45} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF47} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hF48} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hF49} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hF4B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b100, 12'hF4C} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hF4D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hF4E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF4F} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b100, 12'hF51} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF53} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b100, 12'hF55} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hF57} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hF58} : s_CHIP_26B_45133_reg = 8'h93;
         {3'b100, 12'hF59} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hF5B} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hF5D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF5F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b100, 12'hF60} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'hF62} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF63} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hF64} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hF65} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hF66} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF67} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b100, 12'hF68} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hF69} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hF6B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hF6D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF6E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF6F} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hF70} : s_CHIP_26B_45133_reg = 8'h23;
         {3'b100, 12'hF72} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF73} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hF75} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF76} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF77} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hF79} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF7B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b100, 12'hF7D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hF7F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b100, 12'hF80} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hF81} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hF83} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hF84} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hF87} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b100, 12'hF88} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hF8B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hF8C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b100, 12'hF8D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hF8F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hF90} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hF91} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hF93} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b100, 12'hF94} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'hF95} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hF96} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hF97} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b100, 12'hF98} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b100, 12'hF99} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b100, 12'hF9A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hF9B} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b100, 12'hF9C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hF9D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hF9E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hF9F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b100, 12'hFA0} : s_CHIP_26B_45133_reg = 8'hB3;
         {3'b100, 12'hFA1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hFA2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hFA3} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b100, 12'hFA5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hFA7} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hFA8} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b100, 12'hFA9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hFAA} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hFAB} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b100, 12'hFAC} : s_CHIP_26B_45133_reg = 8'hE4;
         {3'b100, 12'hFAD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFAE} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hFAF} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hFB0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFB1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFB3} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b100, 12'hFB4} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hFB5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hFB6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hFB7} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hFB8} : s_CHIP_26B_45133_reg = 8'hA3;
         {3'b100, 12'hFB9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFBB} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hFBD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hFBE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFBF} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b100, 12'hFC1} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hFC2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFC3} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b100, 12'hFC4} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hFC5} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'hFC6} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b100, 12'hFC7} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b100, 12'hFC9} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b100, 12'hFCA} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFCB} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b100, 12'hFCC} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hFCD} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b100, 12'hFCE} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b100, 12'hFCF} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b100, 12'hFD0} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b100, 12'hFD1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hFD3} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hFD5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hFD6} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hFD7} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b100, 12'hFD8} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b100, 12'hFD9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFDA} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hFDB} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b100, 12'hFDC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFDD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b100, 12'hFDE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hFDF} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b100, 12'hFE0} : s_CHIP_26B_45133_reg = 8'h03;
         {3'b100, 12'hFE3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b100, 12'hFE4} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b100, 12'hFE5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hFE7} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b100, 12'hFE8} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b100, 12'hFE9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hFEA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b100, 12'hFEB} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b100, 12'hFEC} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hFED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hFEF} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b100, 12'hFF0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b100, 12'hFF1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hFF2} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b100, 12'hFF3} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b100, 12'hFF4} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b100, 12'hFF5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b100, 12'hFF7} : s_CHIP_26B_45133_reg = 8'h6C;
         {3'b100, 12'hFF9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b100, 12'hFFB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b100, 12'hFFD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b100, 12'hFFF} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h000} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h001} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h003} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b101, 12'h005} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h007} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b101, 12'h008} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h009} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h00B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h00C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b101, 12'h00D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h00E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h00F} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b101, 12'h010} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h011} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h012} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h013} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h014} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h015} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h017} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h018} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h019} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h01B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h01C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h01D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h01F} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b101, 12'h020} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h021} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h023} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h024} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h025} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h027} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h028} : s_CHIP_26B_45133_reg = 8'h7F;
         {3'b101, 12'h029} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h02B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h02D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h02F} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b101, 12'h030} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h031} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h033} : s_CHIP_26B_45133_reg = 8'h38;
         {3'b101, 12'h034} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h035} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h037} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h038} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h039} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h03B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h03C} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b101, 12'h03F} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b101, 12'h040} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b101, 12'h041} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h043} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h044} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b101, 12'h045} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h047} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b101, 12'h049} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h04B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h04D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h04F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h051} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h053} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b101, 12'h055} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b101, 12'h057} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h058} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h059} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b101, 12'h05B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h05C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b101, 12'h05D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h05F} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h060} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h061} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h063} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h064} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b101, 12'h065} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h067} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h068} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h069} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h06B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h06C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h06D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h06F} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h070} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h071} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h073} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h074} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h075} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h077} : s_CHIP_26B_45133_reg = 8'h37;
         {3'b101, 12'h078} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b101, 12'h079} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h07B} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b101, 12'h07D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h07F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h080} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h081} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h083} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b101, 12'h084} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h085} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h086} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h087} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b101, 12'h088} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h089} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h08B} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b101, 12'h08C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h08D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h08F} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h090} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b101, 12'h091} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h092} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h093} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h094} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h095} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h096} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h097} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h098} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h099} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h09B} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h09C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h09D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h09F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h0A0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h0A1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h0A2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h0A3} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b101, 12'h0A5} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b101, 12'h0A6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h0A7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h0A8} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h0A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h0AB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h0AC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h0AD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h0AE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h0AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h0B0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h0B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h0B3} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b101, 12'h0B5} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b101, 12'h0B7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h0B9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b101, 12'h0BB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h0BC} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h0BD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h0BF} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h0C0} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b101, 12'h0C1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h0C2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h0C3} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h0C4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h0C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h0C7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h0C9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h0CA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h0CB} : s_CHIP_26B_45133_reg = 8'h37;
         {3'b101, 12'h0CC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h0CD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h0CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h0D0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h0D2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h0D3} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b101, 12'h0D4} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h0D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h0D7} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b101, 12'h0D8} : s_CHIP_26B_45133_reg = 8'h15;
         {3'b101, 12'h0DA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h0DB} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b101, 12'h0DC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b101, 12'h0DD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h0DF} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h0E0} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h0E2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h0E3} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b101, 12'h0E4} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b101, 12'h0E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h0E7} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h0E8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h0E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h0EA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h0EB} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b101, 12'h0EC} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h0ED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h0EF} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h0F0} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b101, 12'h0F1} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h0F2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h0F3} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h0F4} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h0F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h0F7} : s_CHIP_26B_45133_reg = 8'h66;
         {3'b101, 12'h0F8} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h0F9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h0FB} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h0FC} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b101, 12'h0FD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h0FF} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b101, 12'h100} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h101} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h103} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h104} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b101, 12'h105} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h107} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h108} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b101, 12'h109} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h10A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h10B} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b101, 12'h10C} : s_CHIP_26B_45133_reg = 8'hD4;
         {3'b101, 12'h10D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h10F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h110} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b101, 12'h111} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h113} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b101, 12'h114} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h115} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h117} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b101, 12'h119} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h11A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h11B} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b101, 12'h11C} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b101, 12'h11D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h11E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h11F} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h120} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b101, 12'h121} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h123} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h124} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b101, 12'h126} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h127} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b101, 12'h128} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h129} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h12B} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h12C} : s_CHIP_26B_45133_reg = 8'h44;
         {3'b101, 12'h12D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h12E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h12F} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h130} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b101, 12'h131} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h133} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h134} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h135} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h137} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h138} : s_CHIP_26B_45133_reg = 8'hF4;
         {3'b101, 12'h139} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h13B} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b101, 12'h13C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b101, 12'h13D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h13E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h13F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h140} : s_CHIP_26B_45133_reg = 8'hE4;
         {3'b101, 12'h141} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h143} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h144} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h147} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b101, 12'h148} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h149} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h14B} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b101, 12'h14D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h14F} : s_CHIP_26B_45133_reg = 8'h77;
         {3'b101, 12'h150} : s_CHIP_26B_45133_reg = 8'h15;
         {3'b101, 12'h153} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b101, 12'h155} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h157} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b101, 12'h158} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h159} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h15B} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b101, 12'h15C} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h15D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h15F} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b101, 12'h160} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h161} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h163} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h165} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h166} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h167} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b101, 12'h168} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h169} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h16B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h16C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h16D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h16F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h170} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b101, 12'h171} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h173} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h174} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h175} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h177} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h178} : s_CHIP_26B_45133_reg = 8'hE4;
         {3'b101, 12'h17B} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b101, 12'h17C} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h17D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h17F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h180} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b101, 12'h183} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h184} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b101, 12'h185} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b101, 12'h186} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h187} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h189} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h18B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h18C} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b101, 12'h18D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h18F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h190} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h191} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h192} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h193} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h195} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h197} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b101, 12'h198} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h199} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h19A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h19B} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h19C} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b101, 12'h19D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h19F} : s_CHIP_26B_45133_reg = 8'h59;
         {3'b101, 12'h1A1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h1A2} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h1A3} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h1A4} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b101, 12'h1A5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h1A7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h1A8} : s_CHIP_26B_45133_reg = 8'hFF;
         {3'b101, 12'h1A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1AB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h1AD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1AF} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b101, 12'h1B0} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b101, 12'h1B1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1B3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h1B5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h1B6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h1B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h1B8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h1B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1BB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h1BC} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h1BD} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h1BF} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h1C0} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b101, 12'h1C1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h1C3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h1C4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h1C5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1C6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h1C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h1C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1CB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b101, 12'h1CC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h1CF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h1D0} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h1D2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h1D3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h1D5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1D7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h1D8} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h1D9} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h1DB} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h1DC} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h1DD} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h1DE} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h1DF} : s_CHIP_26B_45133_reg = 8'h02;
         {3'b101, 12'h1E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1E3} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h1E5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h1E6} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h1E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h1E8} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b101, 12'h1E9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h1EA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h1EB} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b101, 12'h1EC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h1ED} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b101, 12'h1EF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h1F0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h1F1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h1F3} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h1F4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h1F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1F7} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h1F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1FB} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h1FC} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h1FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h1FF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h200} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h201} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h202} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h203} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h204} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h205} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h206} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h207} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h208} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h209} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h20B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h20D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h20F} : s_CHIP_26B_45133_reg = 8'h73;
         {3'b101, 12'h211} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h212} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h213} : s_CHIP_26B_45133_reg = 8'h17;
         {3'b101, 12'h214} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h216} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h217} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b101, 12'h219} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h21A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h21B} : s_CHIP_26B_45133_reg = 8'h72;
         {3'b101, 12'h21C} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b101, 12'h21D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h21F} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b101, 12'h221} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h222} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h223} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b101, 12'h224} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h225} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h227} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h228} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h229} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h22B} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h22C} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h22D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h22E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h22F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h230} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h231} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h233} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h234} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h236} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h237} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b101, 12'h238} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h239} : s_CHIP_26B_45133_reg = 8'hB4;
         {3'b101, 12'h23A} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h23B} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b101, 12'h23C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h23D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h23F} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h240} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h241} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h243} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h244} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h245} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h247} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h249} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h24B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h24C} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h24D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h24F} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b101, 12'h250} : s_CHIP_26B_45133_reg = 8'h15;
         {3'b101, 12'h252} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h253} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b101, 12'h254} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b101, 12'h255} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h257} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b101, 12'h258} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h259} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h25B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h25C} : s_CHIP_26B_45133_reg = 8'h24;
         {3'b101, 12'h25D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h25E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h25F} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h260} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h261} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h262} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h263} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h265} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h266} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h267} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b101, 12'h268} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h269} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h26A} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h26B} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b101, 12'h26D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h26E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h26F} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h270} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h271} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h273} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h274} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h275} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h277} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b101, 12'h278} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h279} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h27B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h27D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h27F} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b101, 12'h280} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b101, 12'h281} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h283} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b101, 12'h284} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h285} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h287} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h288} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h289} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h28B} : s_CHIP_26B_45133_reg = 8'h25;
         {3'b101, 12'h28C} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h28D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h28F} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h290} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h291} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h293} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h294} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h295} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b101, 12'h297} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h298} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h299} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b101, 12'h29A} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b101, 12'h29B} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b101, 12'h29D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h29E} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h29F} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b101, 12'h2A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h2A3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h2A5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h2A6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h2A7} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b101, 12'h2A8} : s_CHIP_26B_45133_reg = 8'hA5;
         {3'b101, 12'h2A9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h2AB} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b101, 12'h2AC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h2AD} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h2AF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h2B0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b101, 12'h2B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h2B3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h2B4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h2B5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h2B7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h2B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h2BB} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b101, 12'h2BC} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h2BE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h2BF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h2C0} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h2C1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h2C2} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h2C3} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h2C4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h2C5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h2C7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h2C9} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b101, 12'h2CB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h2CD} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b101, 12'h2CF} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b101, 12'h2D1} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b101, 12'h2D3} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h2D4} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h2D5} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b101, 12'h2D6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h2D7} : s_CHIP_26B_45133_reg = 8'h63;
         {3'b101, 12'h2D8} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b101, 12'h2D9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h2DB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h2DC} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h2DD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h2DE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h2DF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h2E0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h2E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h2E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h2E5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h2E6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h2E7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h2E9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h2EB} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h2ED} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h2EF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h2F1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h2F3} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h2F4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h2F5} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h2F7} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b101, 12'h2F9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h2FB} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b101, 12'h2FC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h2FF} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b101, 12'h301} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h303} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b101, 12'h304} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h305} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h307} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h309} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h30B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h30D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h30E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h30F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b101, 12'h311} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h313} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h314} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b101, 12'h315} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h316} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h317} : s_CHIP_26B_45133_reg = 8'h2A;
         {3'b101, 12'h318} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h319} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b101, 12'h31B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h31C} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b101, 12'h31D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h31E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h31F} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b101, 12'h320} : s_CHIP_26B_45133_reg = 8'hB4;
         {3'b101, 12'h321} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h323} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h324} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b101, 12'h325} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h327} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b101, 12'h329} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b101, 12'h32A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h32B} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b101, 12'h32C} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h32D} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h32E} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h32F} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b101, 12'h331} : s_CHIP_26B_45133_reg = 8'hB1;
         {3'b101, 12'h332} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h333} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b101, 12'h335} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b101, 12'h336} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h337} : s_CHIP_26B_45133_reg = 8'hB9;
         {3'b101, 12'h339} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h33A} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h33B} : s_CHIP_26B_45133_reg = 8'hF9;
         {3'b101, 12'h33C} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h33D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h33F} : s_CHIP_26B_45133_reg = 8'h1A;
         {3'b101, 12'h340} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b101, 12'h341} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h342} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h343} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h344} : s_CHIP_26B_45133_reg = 8'hA4;
         {3'b101, 12'h345} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h347} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b101, 12'h348} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h349} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h34B} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b101, 12'h34C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b101, 12'h34D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h34F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h351} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h352} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h353} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b101, 12'h354} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h355} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h357} : s_CHIP_26B_45133_reg = 8'h71;
         {3'b101, 12'h358} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h359} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h35B} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h35C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h35D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h35F} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b101, 12'h360} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h361} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h363} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b101, 12'h364} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h365} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h367} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h369} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h36B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h36D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h36F} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b101, 12'h371} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h372} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h373} : s_CHIP_26B_45133_reg = 8'h27;
         {3'b101, 12'h374} : s_CHIP_26B_45133_reg = 8'h15;
         {3'b101, 12'h375} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h376} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h377} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h379} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h37B} : s_CHIP_26B_45133_reg = 8'h6F;
         {3'b101, 12'h37D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h37F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h380} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h381} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h383} : s_CHIP_26B_45133_reg = 8'h51;
         {3'b101, 12'h385} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h387} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h388} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h389} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h38B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h38C} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h38F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h391} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h393} : s_CHIP_26B_45133_reg = 8'h11;
         {3'b101, 12'h395} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b101, 12'h397} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b101, 12'h398} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h39A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h39B} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h39D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h39E} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h39F} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b101, 12'h3A0} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b101, 12'h3A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h3A3} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h3A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h3A7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h3A8} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b101, 12'h3A9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h3AA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h3AB} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b101, 12'h3AC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h3AD} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h3AF} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h3B0} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h3B1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h3B3} : s_CHIP_26B_45133_reg = 8'h34;
         {3'b101, 12'h3B4} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h3B5} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h3B7} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h3B8} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h3B9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h3BB} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h3BC} : s_CHIP_26B_45133_reg = 8'hD4;
         {3'b101, 12'h3BF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h3C1} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h3C2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h3C3} : s_CHIP_26B_45133_reg = 8'h61;
         {3'b101, 12'h3C4} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h3C5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h3C7} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h3C8} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h3C9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h3CB} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h3CC} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h3CD} : s_CHIP_26B_45133_reg = 8'h14;
         {3'b101, 12'h3CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h3D0} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h3D1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h3D3} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b101, 12'h3D4} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b101, 12'h3D7} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h3D8} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h3D9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h3DB} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h3DC} : s_CHIP_26B_45133_reg = 8'h75;
         {3'b101, 12'h3DD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h3DF} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h3E0} : s_CHIP_26B_45133_reg = 8'hC0;
         {3'b101, 12'h3E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h3E3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h3E4} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h3E5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h3E7} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h3E8} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b101, 12'h3E9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h3EB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h3EC} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h3ED} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h3EF} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h3F0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h3F1} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h3F3} : s_CHIP_26B_45133_reg = 8'h79;
         {3'b101, 12'h3F4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h3F5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h3F7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h3F8} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h3F9} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h3FB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h3FC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h3FD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h3FF} : s_CHIP_26B_45133_reg = 8'h7B;
         {3'b101, 12'h400} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h401} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h402} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h403} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b101, 12'h405} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h407} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h408} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h409} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h40B} : s_CHIP_26B_45133_reg = 8'h16;
         {3'b101, 12'h40C} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h40D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h40F} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b101, 12'h410} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h411} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h412} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h413} : s_CHIP_26B_45133_reg = 8'h22;
         {3'b101, 12'h414} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b101, 12'h415} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h417} : s_CHIP_26B_45133_reg = 8'h7A;
         {3'b101, 12'h418} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h41B} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h41D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h41F} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h421} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h422} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h423} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h424} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h425} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h426} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h427} : s_CHIP_26B_45133_reg = 8'h13;
         {3'b101, 12'h429} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h42B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h42C} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h42D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h42F} : s_CHIP_26B_45133_reg = 8'h12;
         {3'b101, 12'h430} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h431} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h433} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h434} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h436} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h437} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h438} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h439} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h43B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h43C} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b101, 12'h43D} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h43F} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b101, 12'h440} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h441} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h443} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h444} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h445} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h447} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h448} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b101, 12'h449} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h44B} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h44C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h44D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h44F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h450} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h452} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h453} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h455} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h457} : s_CHIP_26B_45133_reg = 8'h1D;
         {3'b101, 12'h458} : s_CHIP_26B_45133_reg = 8'hB0;
         {3'b101, 12'h459} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h45A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h45B} : s_CHIP_26B_45133_reg = 8'h32;
         {3'b101, 12'h45C} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b101, 12'h45D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h45F} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h460} : s_CHIP_26B_45133_reg = 8'h25;
         {3'b101, 12'h463} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h464} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h465} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b101, 12'h467} : s_CHIP_26B_45133_reg = 8'h31;
         {3'b101, 12'h468} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h469} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h46B} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h46C} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h46D} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h46F} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h470} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h471} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h473} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h474} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h475} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h476} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h477} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h478} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h479} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h47A} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h47B} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h47C} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h47D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h47F} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h481} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h483} : s_CHIP_26B_45133_reg = 8'h33;
         {3'b101, 12'h484} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h485} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h487} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h488} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h489} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h48B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h48C} : s_CHIP_26B_45133_reg = 8'h85;
         {3'b101, 12'h48D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h48F} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h491} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h493} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h495} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h497} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h498} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h499} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h49B} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b101, 12'h49D} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h49F} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h4A0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h4A1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h4A3} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b101, 12'h4A4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h4A5} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h4A7} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h4A8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b101, 12'h4A9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h4AA} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h4AB} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h4AD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h4AE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h4AF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h4B1} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h4B3} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h4B4} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h4B5} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h4B7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h4B8} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h4B9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h4BB} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b101, 12'h4BD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h4BF} : s_CHIP_26B_45133_reg = 8'h39;
         {3'b101, 12'h4C0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b101, 12'h4C1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h4C2} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h4C3} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b101, 12'h4C5} : s_CHIP_26B_45133_reg = 8'h54;
         {3'b101, 12'h4C6} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h4C7} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h4C8} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b101, 12'h4C9} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h4CB} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h4CD} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h4CE} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h4CF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h4D0} : s_CHIP_26B_45133_reg = 8'hE0;
         {3'b101, 12'h4D1} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h4D3} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b101, 12'h4D5} : s_CHIP_26B_45133_reg = 8'h94;
         {3'b101, 12'h4D7} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h4D9} : s_CHIP_26B_45133_reg = 8'h50;
         {3'b101, 12'h4DB} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h4DD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h4DE} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h4DF} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h4E0} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b101, 12'h4E1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h4E3} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b101, 12'h4E4} : s_CHIP_26B_45133_reg = 8'hA0;
         {3'b101, 12'h4E5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h4E6} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h4E7} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b101, 12'h4E8} : s_CHIP_26B_45133_reg = 8'hF5;
         {3'b101, 12'h4E9} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h4EB} : s_CHIP_26B_45133_reg = 8'h19;
         {3'b101, 12'h4EC} : s_CHIP_26B_45133_reg = 8'h15;
         {3'b101, 12'h4EF} : s_CHIP_26B_45133_reg = 8'h6E;
         {3'b101, 12'h4F0} : s_CHIP_26B_45133_reg = 8'h10;
         {3'b101, 12'h4F1} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h4F3} : s_CHIP_26B_45133_reg = 8'h76;
         {3'b101, 12'h4F4} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h4F5} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h4F7} : s_CHIP_26B_45133_reg = 8'h3B;
         {3'b101, 12'h4F8} : s_CHIP_26B_45133_reg = 8'h45;
         {3'b101, 12'h4F9} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h4FA} : s_CHIP_26B_45133_reg = 8'h01;
         {3'b101, 12'h4FB} : s_CHIP_26B_45133_reg = 8'h6B;
         {3'b101, 12'h4FC} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b101, 12'h4FD} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h500} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h503} : s_CHIP_26B_45133_reg = 8'h65;
         {3'b101, 12'h504} : s_CHIP_26B_45133_reg = 8'h70;
         {3'b101, 12'h505} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h507} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h508} : s_CHIP_26B_45133_reg = 8'hF0;
         {3'b101, 12'h509} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h50B} : s_CHIP_26B_45133_reg = 8'h74;
         {3'b101, 12'h50C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h50D} : s_CHIP_26B_45133_reg = 8'h30;
         {3'b101, 12'h50F} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h510} : s_CHIP_26B_45133_reg = 8'h90;
         {3'b101, 12'h511} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h512} : s_CHIP_26B_45133_reg = 8'h40;
         {3'b101, 12'h513} : s_CHIP_26B_45133_reg = 8'h28;
         {3'b101, 12'h514} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h515} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h517} : s_CHIP_26B_45133_reg = 8'h1B;
         {3'b101, 12'h518} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h519} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h51B} : s_CHIP_26B_45133_reg = 8'h3A;
         {3'b101, 12'h51C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h51D} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h51F} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h520} : s_CHIP_26B_45133_reg = 8'hD0;
         {3'b101, 12'h521} : s_CHIP_26B_45133_reg = 8'h81;
         {3'b101, 12'h522} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h523} : s_CHIP_26B_45133_reg = 8'h26;
         {3'b101, 12'h524} : s_CHIP_26B_45133_reg = 8'h04;
         {3'b101, 12'h525} : s_CHIP_26B_45133_reg = 8'h84;
         {3'b101, 12'h527} : s_CHIP_26B_45133_reg = 8'h20;
         {3'b101, 12'h528} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h529} : s_CHIP_26B_45133_reg = 8'h80;
         {3'b101, 12'h52B} : s_CHIP_26B_45133_reg = 8'h60;
         {3'b101, 12'h52C} : s_CHIP_26B_45133_reg = 8'hB5;
         {3'b101, 12'h52E} : s_CHIP_26B_45133_reg = 8'h41;
         {3'b101, 12'h52F} : s_CHIP_26B_45133_reg = 8'h62;
         {3'b101, 12'h530} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h534} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h538} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h53C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h540} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h544} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h548} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h54C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h550} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h554} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h558} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h55C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h560} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h564} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h568} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h56C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h570} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h574} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h578} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h57C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h580} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h584} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h588} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h58C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h590} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h594} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h598} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h59C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5A0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5A4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5A8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5AC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5B0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5B4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5B8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5BC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5C0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5C4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5C8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5CC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5D0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5D4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5D8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5DC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5E0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5E4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5E8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5EC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5F0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5F4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5F8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h5FC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h600} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h604} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h608} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h60C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h610} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h614} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h618} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h61C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h620} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h624} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h628} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h62C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h630} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h634} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h638} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h63C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h640} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h644} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h648} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h64C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h650} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h654} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h658} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h65C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h660} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h664} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h668} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h66C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h670} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h674} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h678} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h67C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h680} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h684} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h688} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h68C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h690} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h694} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h698} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h69C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6A0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6A4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6A8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6AC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6B0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6B4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6B8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6BC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6C0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6C4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6C8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6CC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6D0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6D4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6D8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6DC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6E0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6E4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6E8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6EC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6F0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6F4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6F8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h6FC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h700} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h704} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h708} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h70C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h710} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h714} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h718} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h71C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h720} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h724} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h728} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h72C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h730} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h734} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h738} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h73C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h740} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h744} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h748} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h74C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h750} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h754} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h758} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h75C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h760} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h764} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h768} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h76C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h770} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h774} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h778} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h77C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h780} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h784} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h788} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h78C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h790} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h794} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h798} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h79C} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7A0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7A4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7A8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7AC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7B0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7B4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7B8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7BC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7C0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7C4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7C8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7CC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7D0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7D4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7D8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7DC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7E0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7E4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7E8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7EC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7F0} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7F4} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7F8} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h7FC} : s_CHIP_26B_45133_reg = 8'h05;
         {3'b101, 12'h800} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h804} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h808} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h80C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h810} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h814} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h818} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h81C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h820} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h824} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h828} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h82C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h830} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h834} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h838} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h83C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h840} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h844} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h848} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h84C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h850} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h854} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h858} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h85C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h860} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h864} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h868} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h86C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h870} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h874} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h878} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h87C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h880} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h884} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h888} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h88C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h890} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h894} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h898} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h89C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8A0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8A4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8A8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8AC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8B0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8B4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8B8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8BC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8C0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8C4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8C8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8CC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8D0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8D4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8D8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8DC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8E0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8E4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8E8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8EC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8F0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8F4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8F8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h8FC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h900} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h904} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h908} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h90C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h910} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h914} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h918} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h91C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h920} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h924} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h928} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h92C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h930} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h934} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h938} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h93C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h940} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h944} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h948} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h94C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h950} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h954} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h958} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h95C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h960} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h964} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h968} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h96C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h970} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h974} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h978} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h97C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h980} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h984} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h988} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h98C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h990} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h994} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h998} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h99C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9A0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9A4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9A8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9AC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9B0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9B4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9B8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9BC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9C0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9C4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9C8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9CC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9D0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9D4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9D8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9DC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9E0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9E4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9E8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9EC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9F0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9F4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9F8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'h9FC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA00} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA04} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA08} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA0C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA10} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA14} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA18} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA1C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA20} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA24} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA28} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA2C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA30} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA34} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA38} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA3C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA40} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA44} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA48} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA4C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA50} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA54} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA58} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA5C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA60} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA64} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA68} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA6C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA70} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA74} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA78} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA7C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA80} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA84} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA88} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA8C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA90} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA94} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA98} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hA9C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAA0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAA4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAA8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAAC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAB0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAB4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAB8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hABC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAC0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAC4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAC8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hACC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAD0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAD4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAD8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hADC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAE0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAE4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAE8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAEC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAF0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAF4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAF8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hAFC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB00} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB04} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB08} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB0C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB10} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB14} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB18} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB1C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB20} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB24} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB28} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB2C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB30} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB34} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB38} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB3C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB40} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB44} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB48} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB4C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB50} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB54} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB58} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB5C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB60} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB64} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB68} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB6C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB70} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB74} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB78} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB7C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB80} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB84} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB88} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB8C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB90} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB94} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB98} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hB9C} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBA0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBA4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBA8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBAC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBB0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBB4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBB8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBBC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBC0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBC4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBC8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBCC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBD0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBD4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBD8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBDC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBE0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBE4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBE8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBEC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBF0} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBF4} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBF8} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hBFC} : s_CHIP_26B_45133_reg = 8'h06;
         {3'b101, 12'hC00} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC04} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC08} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC0C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC10} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC14} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC18} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC1C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC20} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC24} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC28} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC2C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC30} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC34} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC38} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC3C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC40} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC44} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC48} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC4C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC50} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC54} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC58} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC5C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC60} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC64} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC68} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC6C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC70} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC74} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC78} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC7C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC80} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC84} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC88} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC8C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC90} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC94} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC98} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hC9C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCA0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCA4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCA8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCAC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCB0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCB4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCB8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCBC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCC0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCC4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCC8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCCC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCD0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCD4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCD8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCDC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCE0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCE4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCE8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCEC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCF0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCF4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCF8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hCFC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD00} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD04} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD08} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD0C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD10} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD14} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD18} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD1C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD20} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD24} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD28} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD2C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD30} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD34} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD38} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD3C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD40} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD44} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD48} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD4C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD50} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD54} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD58} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD5C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD60} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD64} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD68} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD6C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD70} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD74} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD78} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD7C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD80} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD84} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD88} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD8C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD90} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD94} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD98} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hD9C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDA0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDA4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDA8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDAC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDB0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDB4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDB8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDBC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDC0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDC4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDC8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDCC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDD0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDD4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDD8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDDC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDE0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDE4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDE8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDEC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDF0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDF4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDF8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hDFC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE00} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE04} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE08} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE0C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE10} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE14} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE18} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE1C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE20} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE24} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE28} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE2C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE30} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE34} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE38} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE3C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE40} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE44} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE48} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE4C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE50} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE54} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE58} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE5C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE60} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE64} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE68} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE6C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE70} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE74} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE78} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE7C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE80} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE84} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE88} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE8C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE90} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE94} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE98} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hE9C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEA0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEA4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEA8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEAC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEB0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEB4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEB8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEBC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEC0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEC4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEC8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hECC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hED0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hED4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hED8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEDC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEE0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEE4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEE8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEEC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEF0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEF4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEF8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hEFC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF00} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF04} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF08} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF0C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF10} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF14} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF18} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF1C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF20} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF24} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF28} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF2C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF30} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF34} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF38} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF3C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF40} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF44} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF48} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF4C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF50} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF54} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF58} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF5C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF60} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF64} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF68} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF6C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF70} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF74} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF78} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF7C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF80} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF84} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF88} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF8C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF90} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF94} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF98} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hF9C} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFA0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFA4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFA8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFAC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFB0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFB4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFB8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFBC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFC0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFC4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFC8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFCC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFD0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFD4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFD8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFDC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFE0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFE4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFE8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFEC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFF0} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFF4} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFF8} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b101, 12'hFFC} : s_CHIP_26B_45133_reg = 8'h07;
         {3'b110, 12'h000} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h004} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h008} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h00C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h010} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h014} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h018} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h01C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h020} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h024} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h028} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h02C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h030} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h034} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h038} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h03C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h040} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h044} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h048} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h04C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h050} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h054} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h058} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h05C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h060} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h064} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h068} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h06C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h070} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h074} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h078} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h07C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h080} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h084} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h088} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h08C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h090} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h094} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h098} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h09C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0A0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0A4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0A8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0AC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0B0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0B4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0B8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0BC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0C0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0C4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0C8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0CC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0D0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0D4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0D8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0DC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0E0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0E4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0E8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0EC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0F0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0F4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0F8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h0FC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h100} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h104} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h108} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h10C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h110} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h114} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h118} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h11C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h120} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h124} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h128} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h12C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h130} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h134} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h138} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h13C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h140} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h144} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h148} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h14C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h150} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h154} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h158} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h15C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h160} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h164} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h168} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h16C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h170} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h174} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h178} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h17C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h180} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h184} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h188} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h18C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h190} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h194} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h198} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h19C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1A0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1A4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1A8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1AC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1B0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1B4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1B8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1BC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1C0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1C4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1C8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1CC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1D0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1D4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1D8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1DC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1E0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1E4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1E8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1EC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1F0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1F4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1F8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h1FC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h200} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h204} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h208} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h20C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h210} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h214} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h218} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h21C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h220} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h224} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h228} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h22C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h230} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h234} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h238} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h23C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h240} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h244} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h248} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h24C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h250} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h254} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h258} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h25C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h260} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h264} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h268} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h26C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h270} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h274} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h278} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h27C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h280} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h284} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h288} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h28C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h290} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h294} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h298} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h29C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2A0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2A4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2A8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2AC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2B0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2B4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2B8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2BC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2C0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2C4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2C8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2CC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2D0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2D4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2D8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2DC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2E0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2E4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2E8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2EC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2F0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2F4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2F8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h2FC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h300} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h304} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h308} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h30C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h310} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h314} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h318} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h31C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h320} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h324} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h328} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h32C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h330} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h334} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h338} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h33C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h340} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h344} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h348} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h34C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h350} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h354} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h358} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h35C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h360} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h364} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h368} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h36C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h370} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h374} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h378} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h37C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h380} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h384} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h388} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h38C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h390} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h394} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h398} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h39C} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3A0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3A4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3A8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3AC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3B0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3B4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3B8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3BC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3C0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3C4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3C8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3CC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3D0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3D4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3D8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3DC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3E0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3E4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3E8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3EC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3F0} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3F4} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3F8} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h3FC} : s_CHIP_26B_45133_reg = 8'h08;
         {3'b110, 12'h400} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h404} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h408} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h40C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h410} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h414} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h418} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h41C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h420} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h424} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h428} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h42C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h430} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h434} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h438} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h43C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h440} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h444} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h448} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h44C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h450} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h454} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h458} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h45C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h460} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h464} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h468} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h46C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h470} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h474} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h478} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h47C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h480} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h484} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h488} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h48C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h490} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h494} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h498} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h49C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4A0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4A4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4A8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4AC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4B0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4B4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4B8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4BC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4C0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4C4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4C8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4CC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4D0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4D4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4D8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4DC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4E0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4E4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4E8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4EC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4F0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4F4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4F8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h4FC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h500} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h504} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h508} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h50C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h510} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h514} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h518} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h51C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h520} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h524} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h528} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h52C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h530} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h534} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h538} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h53C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h540} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h544} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h548} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h54C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h550} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h554} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h558} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h55C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h560} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h564} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h568} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h56C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h570} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h574} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h578} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h57C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h580} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h584} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h588} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h58C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h590} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h594} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h598} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h59C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5A0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5A4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5A8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5AC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5B0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5B4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5B8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5BC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5C0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5C4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5C8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5CC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5D0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5D4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5D8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5DC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5E0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5E4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5E8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5EC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5F0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5F4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5F8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h5FC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h600} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h604} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h608} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h60C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h610} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h614} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h618} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h61C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h620} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h624} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h628} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h62C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h630} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h634} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h638} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h63C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h640} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h644} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h648} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h64C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h650} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h654} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h658} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h65C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h660} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h664} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h668} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h66C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h670} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h674} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h678} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h67C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h680} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h684} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h688} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h68C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h690} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h694} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h698} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h69C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6A0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6A4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6A8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6AC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6B0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6B4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6B8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6BC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6C0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6C4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6C8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6CC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6D0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6D4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6D8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6DC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6E0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6E4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6E8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6EC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6F0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6F4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6F8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h6FC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h700} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h704} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h708} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h70C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h710} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h714} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h718} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h71C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h720} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h724} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h728} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h72C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h730} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h734} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h738} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h73C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h740} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h744} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h748} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h74C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h750} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h754} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h758} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h75C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h760} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h764} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h768} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h76C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h770} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h774} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h778} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h77C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h780} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h784} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h788} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h78C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h790} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h794} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h798} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h79C} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7A0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7A4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7A8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7AC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7B0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7B4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7B8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7BC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7C0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7C4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7C8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7CC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7D0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7D4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7D8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7DC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7E0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7E4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7E8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7EC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7F0} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7F4} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7F8} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h7FC} : s_CHIP_26B_45133_reg = 8'h09;
         {3'b110, 12'h800} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h804} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h808} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h80C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h810} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h814} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h818} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h81C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h820} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h824} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h828} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h82C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h830} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h834} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h838} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h83C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h840} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h844} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h848} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h84C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h850} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h854} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h858} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h85C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h860} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h864} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h868} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h86C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h870} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h874} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h878} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h87C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h880} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h884} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h888} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h88C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h890} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h894} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h898} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h89C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8A0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8A4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8A8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8AC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8B0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8B4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8B8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8BC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8C0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8C4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8C8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8CC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8D0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8D4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8D8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8DC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8E0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8E4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8E8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8EC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8F0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8F4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8F8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h8FC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h900} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h904} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h908} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h90C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h910} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h914} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h918} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h91C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h920} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h924} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h928} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h92C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h930} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h934} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h938} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h93C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h940} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h944} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h948} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h94C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h950} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h954} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h958} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h95C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h960} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h964} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h968} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h96C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h970} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h974} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h978} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h97C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h980} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h984} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h988} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h98C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h990} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h994} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h998} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h99C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9A0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9A4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9A8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9AC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9B0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9B4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9B8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9BC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9C0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9C4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9C8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9CC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9D0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9D4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9D8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9DC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9E0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9E4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9E8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9EC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9F0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9F4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9F8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'h9FC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA00} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA04} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA08} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA0C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA10} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA14} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA18} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA1C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA20} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA24} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA28} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA2C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA30} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA34} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA38} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA3C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA40} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA44} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA48} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA4C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA50} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA54} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA58} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA5C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA60} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA64} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA68} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA6C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA70} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA74} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA78} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA7C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA80} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA84} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA88} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA8C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA90} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA94} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA98} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hA9C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAA0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAA4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAA8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAAC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAB0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAB4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAB8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hABC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAC0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAC4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAC8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hACC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAD0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAD4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAD8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hADC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAE0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAE4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAE8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAEC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAF0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAF4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAF8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hAFC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB00} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB04} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB08} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB0C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB10} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB14} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB18} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB1C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB20} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB24} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB28} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB2C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB30} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB34} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB38} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB3C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB40} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB44} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB48} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB4C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB50} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB54} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB58} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB5C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB60} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB64} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB68} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB6C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB70} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB74} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB78} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB7C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB80} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB84} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB88} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB8C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB90} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB94} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB98} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hB9C} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBA0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBA4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBA8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBAC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBB0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBB4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBB8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBBC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBC0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBC4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBC8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBCC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBD0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBD4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBD8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBDC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBE0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBE4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBE8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBEC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBF0} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBF4} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBF8} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hBFC} : s_CHIP_26B_45133_reg = 8'h0A;
         {3'b110, 12'hC00} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC04} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC08} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC0C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC10} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC14} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC18} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC1C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC20} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC24} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC28} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC2C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC30} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC34} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC38} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC3C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC40} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC44} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC48} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC4C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC50} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC54} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC58} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC5C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC60} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC64} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC68} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC6C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC70} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC74} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC78} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC7C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC80} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC84} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC88} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC8C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC90} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC94} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC98} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hC9C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCA0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCA4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCA8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCAC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCB0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCB4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCB8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCBC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCC0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCC4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCC8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCCC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCD0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCD4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCD8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCDC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCE0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCE4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCE8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCEC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCF0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCF4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCF8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hCFC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD00} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD04} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD08} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD0C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD10} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD14} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD18} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD1C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD20} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD24} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD28} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD2C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD30} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD34} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD38} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD3C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD40} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD44} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD48} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD4C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD50} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD54} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD58} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD5C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD60} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD64} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD68} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD6C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD70} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD74} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD78} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD7C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD80} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD84} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD88} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD8C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD90} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD94} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD98} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hD9C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDA0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDA4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDA8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDAC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDB0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDB4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDB8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDBC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDC0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDC4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDC8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDCC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDD0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDD4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDD8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDDC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDE0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDE4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDE8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDEC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDF0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDF4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDF8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hDFC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE00} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE04} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE08} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE0C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE10} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE14} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE18} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE1C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE20} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE24} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE28} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE2C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE30} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE34} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE38} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE3C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE40} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE44} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE48} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE4C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE50} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE54} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE58} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE5C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE60} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE64} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE68} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE6C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE70} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE74} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE78} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE7C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE80} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE84} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE88} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE8C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE90} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE94} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE98} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hE9C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEA0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEA4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEA8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEAC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEB0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEB4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEB8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEBC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEC0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEC4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEC8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hECC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hED0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hED4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hED8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEDC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEE0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEE4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEE8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEEC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEF0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEF4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEF8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hEFC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF00} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF04} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF08} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF0C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF10} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF14} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF18} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF1C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF20} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF24} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF28} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF2C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF30} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF34} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF38} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF3C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF40} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF44} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF48} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF4C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF50} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF54} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF58} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF5C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF60} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF64} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF68} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF6C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF70} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF74} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF78} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF7C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF80} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF84} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF88} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF8C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF90} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF94} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF98} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hF9C} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFA0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFA4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFA8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFAC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFB0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFB4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFB8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFBC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFC0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFC4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFC8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFCC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFD0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFD4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFD8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFDC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFE0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFE4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFE8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFEC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFF0} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFF4} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFF8} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b110, 12'hFFC} : s_CHIP_26B_45133_reg = 8'h0B;
         {3'b111, 12'h000} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h004} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h008} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h00C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h010} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h014} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h018} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h01C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h020} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h024} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h028} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h02C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h030} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h034} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h038} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h03C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h040} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h044} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h048} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h04C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h050} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h054} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h058} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h05C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h060} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h064} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h068} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h06C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h070} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h074} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h078} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h07C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h080} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h084} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h088} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h08C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h090} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h094} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h098} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h09C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0A0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0A4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0A8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0AC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0B0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0B4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0B8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0BC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0C0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0C4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0C8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0CC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0D0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0D4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0D8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0DC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0E0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0E4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0E8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0EC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0F0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0F4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0F8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h0FC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h100} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h104} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h108} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h10C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h110} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h114} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h118} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h11C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h120} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h124} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h128} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h12C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h130} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h134} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h138} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h13C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h140} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h144} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h148} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h14C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h150} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h154} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h158} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h15C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h160} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h164} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h168} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h16C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h170} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h174} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h178} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h17C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h180} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h184} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h188} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h18C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h190} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h194} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h198} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h19C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1A0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1A4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1A8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1AC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1B0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1B4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1B8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1BC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1C0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1C4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1C8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1CC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1D0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1D4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1D8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1DC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1E0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1E4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1E8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1EC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1F0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1F4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1F8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h1FC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h200} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h204} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h208} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h20C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h210} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h214} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h218} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h21C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h220} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h224} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h228} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h22C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h230} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h234} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h238} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h23C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h240} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h244} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h248} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h24C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h250} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h254} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h258} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h25C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h260} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h264} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h268} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h26C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h270} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h274} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h278} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h27C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h280} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h284} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h288} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h28C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h290} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h294} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h298} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h29C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2A0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2A4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2A8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2AC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2B0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2B4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2B8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2BC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2C0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2C4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2C8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2CC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2D0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2D4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2D8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2DC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2E0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2E4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2E8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2EC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2F0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2F4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2F8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h2FC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h300} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h304} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h308} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h30C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h310} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h314} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h318} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h31C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h320} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h324} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h328} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h32C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h330} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h334} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h338} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h33C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h340} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h344} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h348} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h34C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h350} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h354} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h358} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h35C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h360} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h364} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h368} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h36C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h370} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h374} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h378} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h37C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h380} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h384} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h388} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h38C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h390} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h394} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h398} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h39C} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3A0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3A4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3A8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3AC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3B0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3B4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3B8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3BC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3C0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3C4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3C8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3CC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3D0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3D4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3D8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3DC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3E0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3E4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3E8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3EC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3F0} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3F4} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3F8} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h3FC} : s_CHIP_26B_45133_reg = 8'h0C;
         {3'b111, 12'h400} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h404} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h408} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h40C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h410} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h414} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h418} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h41C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h420} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h424} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h428} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h42C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h430} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h434} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h438} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h43C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h440} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h444} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h448} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h44C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h450} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h454} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h458} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h45C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h460} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h464} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h468} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h46C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h470} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h474} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h478} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h47C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h480} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h484} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h488} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h48C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h490} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h494} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h498} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h49C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4A0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4A4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4A8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4AC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4B0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4B4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4B8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4BC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4C0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4C4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4C8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4CC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4D0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4D4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4D8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4DC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4E0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4E4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4E8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4EC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4F0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4F4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4F8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h4FC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h500} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h504} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h508} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h50C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h510} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h514} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h518} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h51C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h520} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h524} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h528} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h52C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h530} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h534} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h538} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h53C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h540} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h544} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h548} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h54C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h550} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h554} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h558} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h55C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h560} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h564} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h568} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h56C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h570} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h574} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h578} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h57C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h580} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h584} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h588} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h58C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h590} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h594} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h598} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h59C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5A0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5A4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5A8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5AC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5B0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5B4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5B8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5BC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5C0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5C4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5C8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5CC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5D0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5D4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5D8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5DC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5E0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5E4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5E8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5EC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5F0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5F4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5F8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h5FC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h600} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h604} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h608} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h60C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h610} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h614} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h618} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h61C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h620} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h624} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h628} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h62C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h630} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h634} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h638} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h63C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h640} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h644} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h648} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h64C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h650} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h654} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h658} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h65C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h660} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h664} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h668} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h66C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h670} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h674} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h678} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h67C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h680} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h684} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h688} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h68C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h690} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h694} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h698} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h69C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6A0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6A4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6A8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6AC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6B0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6B4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6B8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6BC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6C0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6C4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6C8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6CC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6D0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6D4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6D8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6DC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6E0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6E4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6E8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6EC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6F0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6F4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6F8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h6FC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h700} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h704} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h708} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h70C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h710} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h714} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h718} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h71C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h720} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h724} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h728} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h72C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h730} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h734} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h738} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h73C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h740} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h744} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h748} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h74C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h750} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h754} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h758} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h75C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h760} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h764} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h768} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h76C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h770} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h774} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h778} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h77C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h780} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h784} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h788} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h78C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h790} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h794} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h798} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h79C} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7A0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7A4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7A8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7AC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7B0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7B4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7B8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7BC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7C0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7C4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7C8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7CC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7D0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7D4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7D8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7DC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7E0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7E4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7E8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7EC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7F0} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7F4} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7F8} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h7FC} : s_CHIP_26B_45133_reg = 8'h0D;
         {3'b111, 12'h800} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h804} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h808} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h80C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h810} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h814} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h818} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h81C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h820} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h824} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h828} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h82C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h830} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h834} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h838} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h83C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h840} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h844} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h848} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h84C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h850} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h854} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h858} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h85C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h860} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h864} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h868} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h86C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h870} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h874} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h878} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h87C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h880} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h884} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h888} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h88C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h890} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h894} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h898} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h89C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8A0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8A4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8A8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8AC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8B0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8B4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8B8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8BC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8C0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8C4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8C8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8CC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8D0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8D4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8D8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8DC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8E0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8E4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8E8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8EC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8F0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8F4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8F8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h8FC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h900} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h904} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h908} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h90C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h910} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h914} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h918} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h91C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h920} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h924} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h928} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h92C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h930} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h934} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h938} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h93C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h940} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h944} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h948} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h94C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h950} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h954} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h958} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h95C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h960} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h964} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h968} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h96C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h970} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h974} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h978} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h97C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h980} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h984} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h988} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h98C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h990} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h994} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h998} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h99C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9A0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9A4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9A8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9AC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9B0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9B4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9B8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9BC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9C0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9C4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9C8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9CC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9D0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9D4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9D8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9DC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9E0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9E4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9E8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9EC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9F0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9F4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9F8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'h9FC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA00} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA04} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA08} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA0C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA10} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA14} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA18} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA1C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA20} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA24} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA28} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA2C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA30} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA34} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA38} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA3C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA40} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA44} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA48} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA4C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA50} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA54} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA58} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA5C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA60} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA64} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA68} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA6C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA70} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA74} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA78} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA7C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA80} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA84} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA88} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA8C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA90} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA94} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA98} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hA9C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAA0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAA4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAA8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAAC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAB0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAB4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAB8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hABC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAC0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAC4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAC8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hACC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAD0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAD4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAD8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hADC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAE0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAE4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAE8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAEC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAF0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAF4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAF8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hAFC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB00} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB04} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB08} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB0C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB10} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB14} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB18} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB1C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB20} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB24} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB28} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB2C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB30} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB34} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB38} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB3C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB40} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB44} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB48} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB4C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB50} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB54} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB58} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB5C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB60} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB64} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB68} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB6C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB70} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB74} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB78} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB7C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB80} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB84} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB88} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB8C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB90} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB94} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB98} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hB9C} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBA0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBA4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBA8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBAC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBB0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBB4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBB8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBBC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBC0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBC4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBC8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBCC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBD0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBD4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBD8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBDC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBE0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBE4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBE8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBEC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBF0} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBF4} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBF8} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hBFC} : s_CHIP_26B_45133_reg = 8'h0E;
         {3'b111, 12'hC00} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC04} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC08} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC0C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC10} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC14} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC18} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC1C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC20} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC24} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC28} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC2C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC30} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC34} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC38} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC3C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC40} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC44} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC48} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC4C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC50} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC54} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC58} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC5C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC60} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC64} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC68} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC6C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC70} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC74} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC78} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC7C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC80} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC84} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC88} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC8C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC90} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC94} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC98} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hC9C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCA0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCA4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCA8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCAC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCB0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCB4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCB8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCBC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCC0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCC4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCC8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCCC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCD0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCD4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCD8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCDC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCE0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCE4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCE8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCEC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCF0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCF4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCF8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hCFC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD00} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD04} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD08} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD0C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD10} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD14} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD18} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD1C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD20} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD24} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD28} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD2C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD30} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD34} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD38} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD3C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD40} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD44} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD48} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD4C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD50} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD54} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD58} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD5C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD60} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD64} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD68} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD6C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD70} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD74} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD78} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD7C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD80} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD84} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD88} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD8C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD90} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD94} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD98} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hD9C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDA0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDA4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDA8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDAC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDB0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDB4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDB8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDBC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDC0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDC4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDC8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDCC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDD0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDD4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDD8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDDC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDE0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDE4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDE8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDEC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDF0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDF4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDF8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hDFC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE00} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE04} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE08} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE0C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE10} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE14} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE18} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE1C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE20} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE24} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE28} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE2C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE30} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE34} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE38} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE3C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE40} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE44} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE48} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE4C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE50} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE54} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE58} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE5C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE60} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE64} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE68} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE6C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE70} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE74} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE78} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE7C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE80} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE84} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE88} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE8C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE90} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE94} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE98} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hE9C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEA0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEA4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEA8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEAC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEB0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEB4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEB8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEBC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEC0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEC4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEC8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hECC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hED0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hED4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hED8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEDC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEE0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEE4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEE8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEEC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEF0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEF4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEF8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hEFC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF00} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF04} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF08} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF0C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF10} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF14} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF18} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF1C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF20} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF24} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF28} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF2C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF30} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF34} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF38} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF3C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF40} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF44} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF48} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF4C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF50} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF54} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF58} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF5C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF60} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF64} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF68} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF6C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF70} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF74} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF78} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF7C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF80} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF84} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF88} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF8C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF90} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF94} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF98} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hF9C} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFA0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFA4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFA8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFAC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFB0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFB4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFB8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFBC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFC0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFC4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFC8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFCC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFD0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFD4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFD8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFDC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFE0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFE4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFE8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFEC} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFF0} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFF4} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFF8} : s_CHIP_26B_45133_reg = 8'h0F;
         {3'b111, 12'hFFC} : s_CHIP_26B_45133_reg = 8'h0F;
         default : s_CHIP_26B_45133_reg = 8'h00;
      endcase
   end

   assign s_databus[15:8] = s_CHIP_26B_45133_reg;

endmodule
