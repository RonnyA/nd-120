
/**************************************************************************
** ND120 CGA (CPU Gate Array / DELILAH)                                  **
** /CGA/ALU/ARG                                                          **
** ARG REGISTER                                                          **
**                                                                       **
** Page 53                                                               **
** SHEET 1 of 1                                                          **
**                                                                       **
** Last reviewed: 30-JAN-2025                                            **
** Ronny Hansen                                                          **
***************************************************************************/

module CGA_ALU_ARG (
    input        ALUCLK,
    input [15:0] CSBIT_15_0,

    output [15:0] ARG_15_0
);

  /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
  wire [15:0] s_csbits_15_0;
  wire        s_aluclk;

  reg [15:0] regArg;

  /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
  assign s_csbits_15_0[15:0] = CSBIT_15_0;
  assign s_aluclk            = ALUCLK;

  /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign ARG_15_0            = regArg;

  /*******************************************************************************
   ** Here all sub-circuits are defined                                          **
   *******************************************************************************/

  always @(posedge s_aluclk) begin
    regArg <= s_csbits_15_0;
  end


endmodule
