/**************************************************************************
** ND120 Shared                                                          **
**                                                                       **
** Component: MUX81                                                      **
**                                                                       **
** Last reviewed: 9-NOV-2024                                             **
** Ronny Hansen                                                          **
***************************************************************************/

module TTL_74521 (
    input [7:0] A_7_0,
    input [7:0] B_7_0,
    input       E_n,

    output AB_n
);

  /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
  wire [7:0] s_a_7_0;
  wire [7:0] s_b_7_0;
  wire       s_ab_n_out;
  wire       s_e_n;
  wire       s_e;
  wire       s_a_equals_b;

  /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

  /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
  assign s_a_7_0[7:0]  = A_7_0;
  assign s_b_7_0[7:0]  = B_7_0;
  assign s_e_n         = E_n;

  /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
  assign AB_n          = s_ab_n_out;

  /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

  // NOT Gate
  assign s_e = ~s_e_n;

  // Controlled Inverter
  assign s_ab_n_out = (s_e) ? ~s_a_equals_b : 1'b0;

  /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
  Comparator #(
      .nrOfBits(8),
      .twosComplement(1)
  ) ARITH_1 (
      .aEqualsB(s_a_equals_b),
      .aGreaterThanB(),
      .aLessThanB(),
      .dataA(s_a_7_0[7:0]),
      .dataB(s_b_7_0[7:0])
  );


endmodule
