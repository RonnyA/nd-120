/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : IDT6168A_20                                                  **
 **                                                                          **
 *****************************************************************************/

module IDT6168A_20( A_11_0,
                    CE_n,
                    D_3_0,
                    WE_n );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input [11:0] A_11_0;
   input        CE_n;
   input        WE_n;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output [3:0] D_3_0;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire [11:0] s_logisimBus1;
   wire [3:0]  s_logisimBus3;
   wire        s_logisimNet0;
   wire        s_logisimNet2;
   wire        s_logisimNet4;
   wire        s_logisimNet5;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
   assign s_logisimBus1[11:0] = A_11_0;
   assign s_logisimNet4       = CE_n;
   assign s_logisimNet5       = WE_n;

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign D_3_0 = s_logisimBus3[3:0];

   /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

   // NOT Gate
   assign s_logisimNet0 = ~s_logisimNet4;

   // NOT Gate
   assign s_logisimNet2 = ~s_logisimNet5;

endmodule
